
//
// Verific Verilog Description of module adder
//

module adder (clk, rx, tx, jtag_inst1_CAPTURE, jtag_inst1_DRCK, jtag_inst1_RESET, 
            jtag_inst1_RUNTEST, jtag_inst1_SEL, jtag_inst1_SHIFT, jtag_inst1_TCK, 
            jtag_inst1_TDI, jtag_inst1_TMS, jtag_inst1_UPDATE, jtag_inst1_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(2)
    input rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(3)
    output tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(4)
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire tx_2;
    wire n25;
    wire [3:0]n26;
    wire [3:0]b;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(10)
    
    wire add_flag, send;
    wire [3:0]sum;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(11)
    
    wire carry;
    wire [3:0]a;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(10)
    
    wire \uart_rx_inst/r_Rx_Data , \uart_rx_inst/r_Rx_Data_R ;
    wire [8:0]\uart_rx_inst/r_Rx_Byte ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(81)
    wire [2:0]\uart_rx_inst/r_SM_Main ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(88)
    wire [31:0]\uart_rx_inst/r_Clock_Count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(79)
    
    wire rx_ready;
    wire [2:0]\uart_rx_inst/r_Bit_Index ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(80)
    wire [31:0]\uart_tx_inst/r_Clock_Count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(203)
    wire [2:0]\uart_tx_inst/r_Bit_Index ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(204)
    wire [7:0]\uart_tx_inst/r_Tx_Data ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(205)
    wire [2:0]\uart_tx_inst/r_SM_Main ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(211)
    
    wire \edb_top_inst/n2056 , \edb_top_inst/la0/la_run_trig ;
    wire [255:0]\edb_top_inst/la0/la_trig_mask ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3481)
    wire [1:0]\edb_top_inst/la0/la_capture_pattern ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3486)
    wire [1:0]\edb_top_inst/la0/la_trig_pattern ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3474)
    
    wire \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig ;
    wire [63:0]\edb_top_inst/la0/skip_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3476)
    wire [16:0]\edb_top_inst/la0/la_num_trigger ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3489)
    wire [4:0]\edb_top_inst/la0/la_window_depth ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3490)
    
    wire \edb_top_inst/la0/la_soft_reset_in ;
    wire [31:0]\edb_top_inst/la0/address_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3403)
    wire [3:0]\edb_top_inst/la0/opcode ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3402)
    wire [5:0]\edb_top_inst/la0/bit_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3404)
    wire [15:0]\edb_top_inst/la0/word_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3405)
    wire [63:0]\edb_top_inst/la0/data_out_shift_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3400)
    wire [3:0]\edb_top_inst/la0/module_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3460)
    
    wire \edb_top_inst/la0/la_resetn_p1 ;
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    
    wire \edb_top_inst/la0/la_resetn ;
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4254)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4270)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4145)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4238)
    wire [43:0]\edb_top_inst/la0/cap_fifo_din_cu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3472)
    wire [43:0]\edb_top_inst/la0/cap_fifo_din_tu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3472)
    wire [12:0]\edb_top_inst/la0/internal_register_select ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3401)
    wire [16:0]\edb_top_inst/la0/la_trig_pos ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3469)
    wire [31:0]\edb_top_inst/la0/crc_data_out ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3456)
    
    wire \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5650)
    
    wire \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ;
    wire [43:0]\edb_top_inst/la0/genblk4.cap_fifo_din_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4447)
    
    wire \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/tu_trigger ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5867)
    
    wire \edb_top_inst/la0/ts_trigger ;
    wire [3:0]\edb_top_inst/la0/la_biu_inst/curr_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4951)
    
    wire \edb_top_inst/la0/la_biu_inst/run_trig_p2 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top_inst/la0/ts_resetn , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ;
    wire [63:0]\edb_top_inst/la0/data_from_biu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3458)
    wire [1:0]\edb_top_inst/la0/la_biu_inst/axi_fsm_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4949)
    
    wire \edb_top_inst/la0/la_biu_inst/run_trig_p1 , \edb_top_inst/la0/biu_ready ;
    wire [31:0]\edb_top_inst/la0/la_biu_inst/addr_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4990)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5393)
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4654)
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    wire [16:0]\edb_top_inst/la0/la_sample_cnt ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3468)
    wire [44:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4768)
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4983)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4644)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4645)
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ;
    wire [3:0]\edb_top_inst/debug_hub_inst/module_id_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(335)
    wire [81:0]\edb_top_inst/edb_user_dr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(45)
    wire [16:0]\edb_top_inst/la0/n1818 ;
    
    wire \edb_top_inst/la0/add_1054/n2 ;
    wire [31:0]\edb_top_inst/la0/n1837 ;
    
    wire \edb_top_inst/la0/add_98/n2 ;
    wire [5:0]\edb_top_inst/la0/n1984 ;
    
    wire \edb_top_inst/la0/add_1057/n2 ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/n73 ;
    
    wire \edb_top_inst/la0/trigger_skipper_n/add_19/n2 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n124 , \edb_top_inst/la0/trigger_skipper_n/add_19/n122 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n120 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 , \edb_top_inst/la0/trigger_skipper_n/add_19/n118 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n116 , \edb_top_inst/la0/trigger_skipper_n/add_19/n114 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n112 , \edb_top_inst/la0/trigger_skipper_n/add_19/n110 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n108 , \edb_top_inst/la0/trigger_skipper_n/add_19/n106 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n104 , \edb_top_inst/la0/trigger_skipper_n/add_19/n102 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n100 , \edb_top_inst/la0/trigger_skipper_n/add_19/n98 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n96 , \edb_top_inst/la0/trigger_skipper_n/add_19/n94 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n92 , \edb_top_inst/la0/trigger_skipper_n/add_19/n90 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n88 , \edb_top_inst/la0/trigger_skipper_n/add_19/n86 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n84 , \edb_top_inst/la0/trigger_skipper_n/add_19/n82 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n80 , \edb_top_inst/la0/trigger_skipper_n/add_19/n78 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n76 , \edb_top_inst/la0/trigger_skipper_n/add_19/n74 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n72 , \edb_top_inst/la0/trigger_skipper_n/add_19/n70 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n68 , \edb_top_inst/la0/trigger_skipper_n/add_19/n66 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n64 , \edb_top_inst/la0/trigger_skipper_n/add_19/n62 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n60 , \edb_top_inst/la0/trigger_skipper_n/add_19/n58 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n56 , \edb_top_inst/la0/trigger_skipper_n/add_19/n54 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n52 , \edb_top_inst/la0/trigger_skipper_n/add_19/n50 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n48 , \edb_top_inst/la0/trigger_skipper_n/add_19/n46 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n44 , \edb_top_inst/la0/trigger_skipper_n/add_19/n42 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n40 , \edb_top_inst/la0/trigger_skipper_n/add_19/n38 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n36 , \edb_top_inst/la0/trigger_skipper_n/add_19/n34 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n32 , \edb_top_inst/la0/trigger_skipper_n/add_19/n30 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n28 , \edb_top_inst/la0/trigger_skipper_n/add_19/n26 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n24 , \edb_top_inst/la0/trigger_skipper_n/add_19/n22 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n20 , \edb_top_inst/la0/trigger_skipper_n/add_19/n18 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n16 , \edb_top_inst/la0/trigger_skipper_n/add_19/n14 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n12 , \edb_top_inst/la0/trigger_skipper_n/add_19/n10 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n8 , \edb_top_inst/la0/trigger_skipper_n/add_19/n6 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n4 , \edb_top_inst/la0/add_1057/n8 , 
        \edb_top_inst/la0/add_1057/n6 , \edb_top_inst/la0/add_1057/n4 , 
        \edb_top_inst/la0/add_98/n48 , \edb_top_inst/la0/add_98/n46 , \edb_top_inst/la0/add_98/n44 , 
        \edb_top_inst/la0/add_98/n42 , \edb_top_inst/la0/add_98/n40 , \edb_top_inst/la0/add_98/n38 , 
        \edb_top_inst/la0/add_98/n36 , \edb_top_inst/la0/add_98/n34 , \edb_top_inst/la0/add_98/n32 , 
        \edb_top_inst/la0/add_98/n30 , \edb_top_inst/la0/add_98/n28 , \edb_top_inst/la0/add_98/n26 , 
        \edb_top_inst/la0/add_98/n24 , \edb_top_inst/la0/add_98/n22 , \edb_top_inst/la0/add_98/n20 , 
        \edb_top_inst/la0/add_98/n18 , \edb_top_inst/la0/add_98/n16 , \edb_top_inst/la0/add_98/n14 , 
        \edb_top_inst/la0/add_98/n12 , \edb_top_inst/la0/add_98/n10 , \edb_top_inst/la0/add_98/n8 , 
        \edb_top_inst/la0/add_98/n6 , \edb_top_inst/la0/add_98/n4 , \edb_top_inst/la0/add_1054/n16 , 
        \edb_top_inst/la0/add_1054/n14 , \edb_top_inst/la0/add_1054/n12 , 
        \edb_top_inst/la0/add_1054/n10 , \edb_top_inst/la0/add_1054/n8 , 
        \edb_top_inst/la0/add_1054/n6 , \edb_top_inst/la0/add_1054/n4 ;
    wire [44:0]\edb_top_inst/la0/la_biu_inst/fifo_dout ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4959)
    
    wire \edb_top_inst/n2057 , \edb_top_inst/n2058 , \edb_top_inst/n2059 , 
        \edb_top_inst/n2060 , \edb_top_inst/n2061 , \edb_top_inst/n2062 , 
        \edb_top_inst/n2063 , \edb_top_inst/n2064 , \edb_top_inst/n2065 , 
        \edb_top_inst/n2066 , \edb_top_inst/n2067 , \edb_top_inst/n2068 , 
        \edb_top_inst/n2069 , \edb_top_inst/n2070 , \edb_top_inst/n2071 , 
        \edb_top_inst/n2072 , \edb_top_inst/n2073 , \edb_top_inst/n2074 , 
        \edb_top_inst/n2075 , \edb_top_inst/n2076 , \edb_top_inst/n2077 , 
        \edb_top_inst/n2078 , \edb_top_inst/n2079 , \edb_top_inst/n2080 , 
        \edb_top_inst/n2081 , \edb_top_inst/n2082 , \edb_top_inst/n2083 , 
        \edb_top_inst/n2084 , \edb_top_inst/n2085 , \edb_top_inst/n2086 , 
        \edb_top_inst/n2087 , \edb_top_inst/n2088 , \edb_top_inst/n2089 , 
        \edb_top_inst/la0/n619 , \edb_top_inst/la0/n618 , \edb_top_inst/n2090 , 
        \edb_top_inst/n2091 , \edb_top_inst/n2092 , \edb_top_inst/n2093 , 
        \edb_top_inst/n2094 , \edb_top_inst/n2095 , \edb_top_inst/n2096 , 
        \edb_top_inst/n2097 , \edb_top_inst/n2098 ;
    wire [3:0]\edb_top_inst/la0/module_next_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3460)
    
    wire \edb_top_inst/n2099 , \edb_top_inst/n2100 , \edb_top_inst/n2101 , 
        \edb_top_inst/n2102 , \edb_top_inst/n2103 , \edb_top_inst/n2104 , 
        \edb_top_inst/n2105 , \edb_top_inst/n2106 , \edb_top_inst/n2107 , 
        \edb_top_inst/n2108 , \edb_top_inst/n2109 , \edb_top_inst/n2110 , 
        \edb_top_inst/n2111 , \edb_top_inst/n2112 , \edb_top_inst/n2113 , 
        \edb_top_inst/n2114 , \edb_top_inst/n2115 , \edb_top_inst/n2116 , 
        \edb_top_inst/la0/n1022 , \edb_top_inst/n2117 , \edb_top_inst/n2118 , 
        \edb_top_inst/n2119 , \edb_top_inst/n2120 , \edb_top_inst/n2121 , 
        \edb_top_inst/n2122 , \edb_top_inst/la0/regsel_ld_en , \edb_top_inst/n2123 , 
        \edb_top_inst/n2124 , \edb_top_inst/n2125 , \edb_top_inst/la0/n994 , 
        \edb_top_inst/ceg_net2 , \edb_top_inst/n2126 , \edb_top_inst/la0/n1078 , 
        \edb_top_inst/la0/n1023 , \edb_top_inst/la0/n1024 , \edb_top_inst/n2127 , 
        \edb_top_inst/n2128 , \edb_top_inst/la0/n1595 , \edb_top_inst/la0/n1728 , 
        \edb_top_inst/n2129 , \edb_top_inst/la0/n1780 , \edb_top_inst/n2130 , 
        \edb_top_inst/n2131 , \edb_top_inst/n2132 , \edb_top_inst/n2133 , 
        \edb_top_inst/n2134 ;
    wire [31:0]\edb_top_inst/la0/data_to_addr_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3450)
    
    wire \edb_top_inst/n2135 , \edb_top_inst/n2136 , \edb_top_inst/n2137 , 
        \edb_top_inst/n2138 , \edb_top_inst/n2139 , \edb_top_inst/n2140 , 
        \edb_top_inst/n2141 , \edb_top_inst/n2142 , \edb_top_inst/n2143 , 
        \edb_top_inst/n2144 , \edb_top_inst/la0/addr_ct_en , \edb_top_inst/la0/n616 , 
        \edb_top_inst/la0/op_reg_en , \edb_top_inst/n2145 , \edb_top_inst/n2146 , 
        \edb_top_inst/n2147 ;
    wire [5:0]\edb_top_inst/la0/n1998 ;
    
    wire \edb_top_inst/n2148 , \edb_top_inst/n2149 , \edb_top_inst/ceg_net5 ;
    wire [15:0]\edb_top_inst/la0/data_to_word_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3453)
    
    wire \edb_top_inst/n2150 , \edb_top_inst/n2151 , \edb_top_inst/la0/word_ct_en , 
        \edb_top_inst/n2152 , \edb_top_inst/n2153 , \edb_top_inst/n2154 , 
        \edb_top_inst/n2155 , \edb_top_inst/n2156 , \edb_top_inst/n2157 , 
        \edb_top_inst/n2158 , \edb_top_inst/n2159 , \edb_top_inst/n2160 , 
        \edb_top_inst/n2161 , \edb_top_inst/n2162 , \edb_top_inst/n2163 , 
        \edb_top_inst/n2164 , \edb_top_inst/n2165 , \edb_top_inst/n2166 , 
        \edb_top_inst/n2167 , \edb_top_inst/n2168 ;
    wire [63:0]\edb_top_inst/la0/n2217 ;
    
    wire \edb_top_inst/n2169 , \edb_top_inst/ceg_net8 , \edb_top_inst/la0/n2568 , 
        \edb_top_inst/n2170 , \edb_top_inst/n2171 , \edb_top_inst/la0/n2581 , 
        \edb_top_inst/n2172 , \edb_top_inst/n2173 , \edb_top_inst/la0/n3470 , 
        \edb_top_inst/la0/n3485 , \edb_top_inst/n2174 , \edb_top_inst/la0/n3683 , 
        \edb_top_inst/la0/n4311 , \edb_top_inst/n2175 , \edb_top_inst/la0/n5144 , 
        \edb_top_inst/la0/n5977 , \edb_top_inst/la0/n6810 , \edb_top_inst/la0/n7643 , 
        \edb_top_inst/n2176 , \edb_top_inst/n2177 , \edb_top_inst/la0/n8532 , 
        \edb_top_inst/la0/n8547 , \edb_top_inst/la0/n8745 , \edb_top_inst/n2178 , 
        \edb_top_inst/la0/n9429 , \edb_top_inst/la0/n9444 , \edb_top_inst/la0/n9642 , 
        \edb_top_inst/n2179 , \edb_top_inst/la0/n10298 , \edb_top_inst/la0/n10313 , 
        \edb_top_inst/la0/n10511 , \edb_top_inst/n2180 , \edb_top_inst/la0/n11163 , 
        \edb_top_inst/la0/n11178 , \edb_top_inst/la0/n11376 , \edb_top_inst/n2181 , 
        \edb_top_inst/la0/n12028 , \edb_top_inst/la0/n12043 , \edb_top_inst/la0/n12241 , 
        \edb_top_inst/n2182 , \edb_top_inst/la0/n12865 , \edb_top_inst/la0/n13698 , 
        \edb_top_inst/n2183 , \edb_top_inst/n2184 , \edb_top_inst/n2185 , 
        \edb_top_inst/n2186 , \edb_top_inst/n2187 , \edb_top_inst/n2188 , 
        \edb_top_inst/n2189 , \edb_top_inst/n2190 , \edb_top_inst/n2191 , 
        \edb_top_inst/n2192 , \edb_top_inst/n2200 , \edb_top_inst/n2201 , 
        \edb_top_inst/n2202 , \edb_top_inst/n2203 , \edb_top_inst/n2204 , 
        \edb_top_inst/n2205 , \edb_top_inst/n2206 , \edb_top_inst/n2207 , 
        \edb_top_inst/n2208 , \edb_top_inst/n2209 , \edb_top_inst/n2210 , 
        \edb_top_inst/n2211 , \edb_top_inst/n2212 , \edb_top_inst/n2213 , 
        \edb_top_inst/n2214 , \edb_top_inst/n2215 , \edb_top_inst/n2216 , 
        \edb_top_inst/n2217 , \edb_top_inst/n2218 , \edb_top_inst/n2219 , 
        \edb_top_inst/n2220 , \edb_top_inst/n2221 , \edb_top_inst/n2222 , 
        \edb_top_inst/n2223 , \edb_top_inst/n2224 , \edb_top_inst/n2225 , 
        \edb_top_inst/n2226 , \edb_top_inst/n2227 , \edb_top_inst/n2228 , 
        \edb_top_inst/n2229 , \edb_top_inst/n2230 , \edb_top_inst/n2231 , 
        \edb_top_inst/n2232 , \edb_top_inst/n2233 , \edb_top_inst/n2234 , 
        \edb_top_inst/n2235 , \edb_top_inst/n2237 , \edb_top_inst/n2055 , 
        \edb_top_inst/n2238 , \edb_top_inst/n2239 , \edb_top_inst/n2240 , 
        \edb_top_inst/n2241 , \edb_top_inst/n2242 , \edb_top_inst/n2243 , 
        \edb_top_inst/n2244 , \edb_top_inst/n2245 , \edb_top_inst/n2246 , 
        \edb_top_inst/n2247 , \edb_top_inst/n2248 , \edb_top_inst/n2249 , 
        \edb_top_inst/n2250 , \edb_top_inst/n2251 , \edb_top_inst/n2252 , 
        \edb_top_inst/n2253 , \edb_top_inst/n2254 , \edb_top_inst/n2255 , 
        \edb_top_inst/n2256 , \edb_top_inst/n2257 , \edb_top_inst/n2258 , 
        \edb_top_inst/n2259 , \edb_top_inst/n2260 , \edb_top_inst/n2261 , 
        \edb_top_inst/n2262 , \edb_top_inst/n2263 , \edb_top_inst/n2264 , 
        \edb_top_inst/n2265 , \edb_top_inst/n2266 , \edb_top_inst/n2267 , 
        \edb_top_inst/n2268 , \edb_top_inst/n2269 , \edb_top_inst/n2270 , 
        \edb_top_inst/n2271 , \edb_top_inst/n2272 , \edb_top_inst/n2273 , 
        \edb_top_inst/n2274 , \edb_top_inst/n2275 , \edb_top_inst/n2276 , 
        \edb_top_inst/n2277 , \edb_top_inst/n2278 , \edb_top_inst/n2279 , 
        \edb_top_inst/n2280 , \edb_top_inst/n2281 , \edb_top_inst/n2282 , 
        \edb_top_inst/n2283 , \edb_top_inst/n2284 , \edb_top_inst/n2285 , 
        \edb_top_inst/n2286 , \edb_top_inst/n2287 , \edb_top_inst/n2288 , 
        \edb_top_inst/n2289 , \edb_top_inst/n2290 , \edb_top_inst/n2291 , 
        \edb_top_inst/n2292 , \edb_top_inst/n2293 , \edb_top_inst/n2294 , 
        \edb_top_inst/n2295 , \edb_top_inst/n2296 , \edb_top_inst/n2297 , 
        \edb_top_inst/n2298 , \edb_top_inst/n2299 , \edb_top_inst/n2300 , 
        \edb_top_inst/n2301 , \edb_top_inst/n2302 , \edb_top_inst/n2303 , 
        \edb_top_inst/n2304 , \edb_top_inst/n2305 , \edb_top_inst/n2306 , 
        \edb_top_inst/n2307 , \edb_top_inst/n2308 , \edb_top_inst/n2309 , 
        \edb_top_inst/n2310 , \edb_top_inst/n2311 , \edb_top_inst/n2312 , 
        \edb_top_inst/n2313 , \edb_top_inst/n2314 , \edb_top_inst/n2315 , 
        \edb_top_inst/n2316 , \edb_top_inst/n2317 , \edb_top_inst/n2318 , 
        \edb_top_inst/n2319 , \edb_top_inst/n2320 , \edb_top_inst/n2321 , 
        \edb_top_inst/n2322 , \edb_top_inst/n2323 , \edb_top_inst/n2324 , 
        \edb_top_inst/n2325 , \edb_top_inst/n2326 , \edb_top_inst/n2327 , 
        \edb_top_inst/n2328 , \edb_top_inst/n2329 , \edb_top_inst/n2330 , 
        \edb_top_inst/n2331 , \edb_top_inst/n2332 , \edb_top_inst/n2333 , 
        \edb_top_inst/n2334 , \edb_top_inst/n2335 , \edb_top_inst/n2336 , 
        \edb_top_inst/n2337 , \edb_top_inst/n2338 , \edb_top_inst/n2339 , 
        \edb_top_inst/n2340 , \edb_top_inst/n2341 , \edb_top_inst/n2342 , 
        \edb_top_inst/n2343 , \edb_top_inst/n2344 , \edb_top_inst/n2345 , 
        \edb_top_inst/n2346 , \edb_top_inst/n2347 , \edb_top_inst/n2348 , 
        \edb_top_inst/n2349 , \edb_top_inst/n2350 , \edb_top_inst/n2351 , 
        \edb_top_inst/n2352 , \edb_top_inst/n2353 , \edb_top_inst/n2354 , 
        \edb_top_inst/n2355 , \edb_top_inst/n2356 , \edb_top_inst/n2357 , 
        \edb_top_inst/n2358 , \edb_top_inst/n2359 , \edb_top_inst/n2360 , 
        \edb_top_inst/n2361 , \edb_top_inst/n2362 , \edb_top_inst/n2363 , 
        \edb_top_inst/n2364 , \edb_top_inst/n2365 , \edb_top_inst/n2366 , 
        \edb_top_inst/n2367 , \edb_top_inst/n2368 , \edb_top_inst/n2369 , 
        \edb_top_inst/n2370 , \edb_top_inst/n2371 , \edb_top_inst/n2372 , 
        \edb_top_inst/n2373 , \edb_top_inst/n2374 , \edb_top_inst/n2375 , 
        \edb_top_inst/n2376 , \edb_top_inst/n2377 , \edb_top_inst/n2378 , 
        \edb_top_inst/n2379 , \edb_top_inst/n2380 , \edb_top_inst/n2381 , 
        \edb_top_inst/n2382 , \edb_top_inst/n2383 , \edb_top_inst/n2384 , 
        \edb_top_inst/n2385 , \edb_top_inst/n2386 , \edb_top_inst/n2387 , 
        \edb_top_inst/n2388 , \edb_top_inst/n2389 , \edb_top_inst/n2390 , 
        \edb_top_inst/n2391 , \edb_top_inst/n2392 , \edb_top_inst/n2393 , 
        \edb_top_inst/n2394 ;
    wire [31:0]\edb_top_inst/la0/axi_crc_i/n118 ;
    
    wire \edb_top_inst/ceg_net11 , \edb_top_inst/n2395 , \edb_top_inst/n2396 , 
        \edb_top_inst/n2397 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2398 , \edb_top_inst/n2399 , \edb_top_inst/n2400 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 ;
    
    wire \edb_top_inst/n2401 , \edb_top_inst/n2402 , \edb_top_inst/n2403 , 
        \edb_top_inst/n2404 , \edb_top_inst/n2405 , \edb_top_inst/n2406 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/n2407 , 
        \edb_top_inst/n2408 , \edb_top_inst/n2409 , \edb_top_inst/n2410 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/n2411 , \edb_top_inst/n2412 , \edb_top_inst/n2413 , 
        \edb_top_inst/n2414 , \edb_top_inst/n2415 , \edb_top_inst/n2416 , 
        \edb_top_inst/n2417 , \edb_top_inst/n2418 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2419 , \edb_top_inst/n2420 , \edb_top_inst/n2421 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2422 , \edb_top_inst/n2423 , \edb_top_inst/n2424 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2425 , \edb_top_inst/n2426 , \edb_top_inst/n2427 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n2428 , 
        \edb_top_inst/n2429 , \edb_top_inst/n2430 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2431 , \edb_top_inst/n2432 , \edb_top_inst/n2433 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 ;
    
    wire \edb_top_inst/n2434 , \edb_top_inst/n2435 , \edb_top_inst/n2436 , 
        \edb_top_inst/n2437 , \edb_top_inst/n2438 , \edb_top_inst/n2439 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/n2440 , 
        \edb_top_inst/n2441 , \edb_top_inst/n2442 , \edb_top_inst/n2443 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/n2444 , \edb_top_inst/n2445 , \edb_top_inst/n2446 , 
        \edb_top_inst/n2447 , \edb_top_inst/n2448 , \edb_top_inst/n2449 , 
        \edb_top_inst/n2450 , \edb_top_inst/n2451 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 ;
    
    wire \edb_top_inst/n2452 , \edb_top_inst/n2453 , \edb_top_inst/n2454 , 
        \edb_top_inst/n2455 , \edb_top_inst/n2456 , \edb_top_inst/n2457 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/n2458 , 
        \edb_top_inst/n2459 , \edb_top_inst/n2460 , \edb_top_inst/n2461 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/n2462 , \edb_top_inst/n2463 , \edb_top_inst/n2464 , 
        \edb_top_inst/n2465 , \edb_top_inst/n2466 , \edb_top_inst/n2467 , 
        \edb_top_inst/n2468 , \edb_top_inst/n2469 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 ;
    
    wire \edb_top_inst/n2470 , \edb_top_inst/n2471 , \edb_top_inst/n2472 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n25 , \edb_top_inst/n2473 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n7 , 
        \edb_top_inst/n2474 , \edb_top_inst/n2475 , \edb_top_inst/n2476 , 
        \edb_top_inst/n2477 , \edb_top_inst/n2478 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 ;
    
    wire \edb_top_inst/n2479 , \edb_top_inst/n2480 , \edb_top_inst/n2481 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n25 , \edb_top_inst/n2482 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/equal_9/n7 , 
        \edb_top_inst/n2483 , \edb_top_inst/n2484 , \edb_top_inst/n2485 , 
        \edb_top_inst/n2486 , \edb_top_inst/n2487 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n34 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 ;
    wire [3:0]\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 ;
    
    wire \edb_top_inst/n2488 , \edb_top_inst/n2490 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n25 , 
        \edb_top_inst/n2491 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/equal_9/n7 , 
        \edb_top_inst/n2492 , \edb_top_inst/n2493 , \edb_top_inst/n2494 , 
        \edb_top_inst/n2495 , \edb_top_inst/n2496 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2497 , \edb_top_inst/n2498 , \edb_top_inst/n2499 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n2500 , \edb_top_inst/n2501 , \edb_top_inst/n2502 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n2503 , 
        \edb_top_inst/n2504 , \edb_top_inst/n2505 , \edb_top_inst/n2506 , 
        \edb_top_inst/n2507 , \edb_top_inst/n2508 , \edb_top_inst/n2509 , 
        \edb_top_inst/n2510 , \edb_top_inst/n2511 , \edb_top_inst/n2512 , 
        \edb_top_inst/n2513 , \edb_top_inst/n2514 , \edb_top_inst/n2515 , 
        \edb_top_inst/n2516 , \edb_top_inst/n2517 , \edb_top_inst/n2518 , 
        \edb_top_inst/n2519 , \edb_top_inst/n2520 , \edb_top_inst/n2521 , 
        \edb_top_inst/n2522 , \edb_top_inst/n2523 , \edb_top_inst/n2524 , 
        \edb_top_inst/n2525 , \edb_top_inst/la0/trigger_tu/n101 , \edb_top_inst/n2526 , 
        \edb_top_inst/n2527 , \edb_top_inst/n2528 , \edb_top_inst/n2529 , 
        \edb_top_inst/n2530 , \edb_top_inst/n2531 , \edb_top_inst/n2532 , 
        \edb_top_inst/n2533 , \edb_top_inst/n2534 , \edb_top_inst/n2535 , 
        \edb_top_inst/n2536 , \edb_top_inst/n2537 , \edb_top_inst/n2538 , 
        \edb_top_inst/n2539 , \edb_top_inst/n2540 , \edb_top_inst/n2541 , 
        \edb_top_inst/n2542 , \edb_top_inst/n2543 , \edb_top_inst/n2544 , 
        \edb_top_inst/n2545 , \edb_top_inst/n2546 , \edb_top_inst/n2547 , 
        \edb_top_inst/n2548 , \edb_top_inst/n2549 , \edb_top_inst/n2550 , 
        \edb_top_inst/n2551 , \edb_top_inst/n2552 , \edb_top_inst/n2553 , 
        \edb_top_inst/n2554 , \edb_top_inst/n2555 , \edb_top_inst/n2556 , 
        \edb_top_inst/n2557 , \edb_top_inst/n2558 , \edb_top_inst/n2559 , 
        \edb_top_inst/n2560 , \edb_top_inst/n2561 , \edb_top_inst/n2562 , 
        \edb_top_inst/n2563 , \edb_top_inst/n2564 , \edb_top_inst/n2565 , 
        \edb_top_inst/n2566 , \edb_top_inst/n2567 , \edb_top_inst/n2568 , 
        \edb_top_inst/n2569 , \edb_top_inst/n2570 , \edb_top_inst/n2571 , 
        \edb_top_inst/n2572 , \edb_top_inst/n2573 , \edb_top_inst/n2574 , 
        \edb_top_inst/n2575 , \edb_top_inst/n2576 , \edb_top_inst/n2577 , 
        \edb_top_inst/n2578 , \edb_top_inst/n2579 , \edb_top_inst/n2580 , 
        \edb_top_inst/n2581 , \edb_top_inst/n2582 , \edb_top_inst/n2583 , 
        \edb_top_inst/n2584 , \edb_top_inst/n2585 , \edb_top_inst/n2586 , 
        \edb_top_inst/n2587 , \edb_top_inst/n2588 , \edb_top_inst/n2589 , 
        \edb_top_inst/n2590 , \edb_top_inst/n2591 , \edb_top_inst/n2592 , 
        \edb_top_inst/n2593 , \edb_top_inst/n2594 , \edb_top_inst/n2595 , 
        \edb_top_inst/n2596 , \edb_top_inst/n2597 , \edb_top_inst/n2598 , 
        \edb_top_inst/n2599 , \edb_top_inst/n2600 , \edb_top_inst/n2601 , 
        \edb_top_inst/n2602 , \edb_top_inst/n2603 , \edb_top_inst/n2604 , 
        \edb_top_inst/n2605 , \edb_top_inst/n2606 , \edb_top_inst/n2607 , 
        \edb_top_inst/n2608 , \edb_top_inst/n2609 , \edb_top_inst/n2610 , 
        \edb_top_inst/n2611 , \edb_top_inst/n2612 , \edb_top_inst/n2613 , 
        \edb_top_inst/n2614 , \edb_top_inst/n2615 , \edb_top_inst/n2616 , 
        \edb_top_inst/n2617 , \edb_top_inst/n2618 , \edb_top_inst/n2619 , 
        \edb_top_inst/n2620 , \edb_top_inst/n2621 , \edb_top_inst/n2622 , 
        \edb_top_inst/n2623 , \edb_top_inst/n2624 , \edb_top_inst/n2625 , 
        \edb_top_inst/n2626 , \edb_top_inst/n2627 , \edb_top_inst/n2628 , 
        \edb_top_inst/n2629 , \edb_top_inst/n2630 , \edb_top_inst/n2631 , 
        \edb_top_inst/n2632 , \edb_top_inst/n2633 , \edb_top_inst/n2634 , 
        \edb_top_inst/n2635 , \edb_top_inst/n2636 , \edb_top_inst/n2637 , 
        \edb_top_inst/n2638 , \edb_top_inst/n2639 , \edb_top_inst/n2640 , 
        \edb_top_inst/n2641 , \edb_top_inst/n2642 , \edb_top_inst/n2643 , 
        \edb_top_inst/n2644 , \edb_top_inst/n2645 , \edb_top_inst/n2646 , 
        \edb_top_inst/n2647 , \edb_top_inst/n2648 , \edb_top_inst/n2649 , 
        \edb_top_inst/n2650 , \edb_top_inst/n2651 , \edb_top_inst/n2652 , 
        \edb_top_inst/n2653 , \edb_top_inst/n2654 , \edb_top_inst/n2655 , 
        \edb_top_inst/n2656 , \edb_top_inst/n2657 , \edb_top_inst/n2658 , 
        \edb_top_inst/n2659 , \edb_top_inst/n2660 , \edb_top_inst/n2661 , 
        \edb_top_inst/n2662 , \edb_top_inst/n2663 , \edb_top_inst/n2664 , 
        \edb_top_inst/n2665 , \edb_top_inst/n2666 , \edb_top_inst/n2667 , 
        \edb_top_inst/n2668 , \edb_top_inst/n2669 , \edb_top_inst/n2670 , 
        \edb_top_inst/n2671 , \edb_top_inst/n2672 , \edb_top_inst/n2673 , 
        \edb_top_inst/n2674 , \edb_top_inst/n2675 , \edb_top_inst/n2676 , 
        \edb_top_inst/n2677 , \edb_top_inst/n2678 ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/n138 ;
    
    wire \edb_top_inst/la0/trigger_skipper_n/n468 , \edb_top_inst/n2679 , 
        \edb_top_inst/n2680 , \edb_top_inst/n2681 , \edb_top_inst/n2682 , 
        \edb_top_inst/n2683 , \edb_top_inst/n2684 , \edb_top_inst/n2685 , 
        \edb_top_inst/n2686 , \edb_top_inst/n2687 , \edb_top_inst/n2688 , 
        \edb_top_inst/n2689 , \edb_top_inst/n2690 , \edb_top_inst/n2691 , 
        \edb_top_inst/n2692 , \edb_top_inst/n2693 , \edb_top_inst/n2694 , 
        \edb_top_inst/n2695 , \edb_top_inst/n2696 , \edb_top_inst/n2697 , 
        \edb_top_inst/n2698 , \edb_top_inst/n2699 , \edb_top_inst/n2700 , 
        \edb_top_inst/n2701 , \edb_top_inst/n2702 , \edb_top_inst/n2703 , 
        \edb_top_inst/n2704 , \edb_top_inst/n2705 , \edb_top_inst/n2706 , 
        \edb_top_inst/n2707 , \edb_top_inst/n2708 , \edb_top_inst/n2709 , 
        \edb_top_inst/n2710 , \edb_top_inst/n2711 , \edb_top_inst/n2712 , 
        \edb_top_inst/n2713 , \edb_top_inst/n2714 , \edb_top_inst/n2715 , 
        \edb_top_inst/n2716 , \edb_top_inst/n2717 , \edb_top_inst/n2718 , 
        \edb_top_inst/n2719 , \edb_top_inst/n2720 , \edb_top_inst/n2721 , 
        \edb_top_inst/n2722 , \edb_top_inst/n2723 , \edb_top_inst/n2724 , 
        \edb_top_inst/n2725 , \edb_top_inst/n2726 , \edb_top_inst/n2727 , 
        \edb_top_inst/n2728 , \edb_top_inst/n2729 , \edb_top_inst/n2730 , 
        \edb_top_inst/n2731 , \edb_top_inst/n2732 , \edb_top_inst/n2733 , 
        \edb_top_inst/n2734 , \edb_top_inst/n2735 , \edb_top_inst/n2736 , 
        \edb_top_inst/n2737 , \edb_top_inst/n2738 , \edb_top_inst/n2739 , 
        \edb_top_inst/n2740 , \edb_top_inst/n2741 , \edb_top_inst/n2742 , 
        \edb_top_inst/n2743 , \edb_top_inst/n2744 , \edb_top_inst/n2745 , 
        \edb_top_inst/n2746 , \edb_top_inst/n2747 , \edb_top_inst/n2748 , 
        \edb_top_inst/n2749 , \edb_top_inst/n2750 , \edb_top_inst/n2751 , 
        \edb_top_inst/n2752 , \edb_top_inst/n2753 , \edb_top_inst/n2754 , 
        \edb_top_inst/n2755 , \edb_top_inst/n2756 , \edb_top_inst/n2757 , 
        \edb_top_inst/n2758 , \edb_top_inst/n2759 , \edb_top_inst/n2760 , 
        \edb_top_inst/n2761 , \edb_top_inst/n2762 , \edb_top_inst/n2763 , 
        \edb_top_inst/n2764 , \edb_top_inst/n2765 , \edb_top_inst/n2766 , 
        \edb_top_inst/n2767 , \edb_top_inst/n2768 , \edb_top_inst/n2769 , 
        \edb_top_inst/n2770 , \edb_top_inst/n2771 , \edb_top_inst/n2772 , 
        \edb_top_inst/n2773 , \edb_top_inst/n2774 , \edb_top_inst/n2775 , 
        \edb_top_inst/n2776 , \edb_top_inst/n2777 , \edb_top_inst/n2778 , 
        \edb_top_inst/n2779 , \edb_top_inst/n2780 , \edb_top_inst/n2781 , 
        \edb_top_inst/n2782 , \edb_top_inst/n2783 , \edb_top_inst/n2784 , 
        \edb_top_inst/n2785 , \edb_top_inst/n2786 , \edb_top_inst/n2787 , 
        \edb_top_inst/n2788 , \edb_top_inst/n2789 , \edb_top_inst/n2790 , 
        \edb_top_inst/n2791 , \edb_top_inst/n2792 , \edb_top_inst/n2793 , 
        \edb_top_inst/n2794 , \edb_top_inst/n2795 , \edb_top_inst/n2796 , 
        \edb_top_inst/n2797 , \edb_top_inst/n2798 , \edb_top_inst/n2799 , 
        \edb_top_inst/n2800 , \edb_top_inst/n2801 , \edb_top_inst/n2802 ;
    wire [3:0]\edb_top_inst/la0/la_biu_inst/next_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4951)
    
    wire \edb_top_inst/la0/la_biu_inst/n98 , \edb_top_inst/n2803 , \edb_top_inst/la0/la_biu_inst/n370 , 
        \edb_top_inst/la0/la_biu_inst/n1318 , \edb_top_inst/la0/la_biu_inst/n1319 , 
        \edb_top_inst/la0/la_biu_inst/n1902 , \edb_top_inst/n2804 , \edb_top_inst/n2805 , 
        \edb_top_inst/n2806 , \edb_top_inst/n2807 , \edb_top_inst/la0/la_biu_inst/n1284 , 
        \edb_top_inst/la0/n19936 , \edb_top_inst/n2808 , \edb_top_inst/n2809 , 
        \edb_top_inst/n2810 , \edb_top_inst/n2811 , \edb_top_inst/n2812 , 
        \edb_top_inst/n2813 , \edb_top_inst/n2814 , \edb_top_inst/n2815 , 
        \edb_top_inst/n2816 , \edb_top_inst/n2817 , \edb_top_inst/n2818 , 
        \edb_top_inst/n2819 , \edb_top_inst/n2820 , \edb_top_inst/n2821 , 
        \edb_top_inst/n2822 , \edb_top_inst/ceg_net18 ;
    wire [1:0]\edb_top_inst/la0/la_biu_inst/next_fsm_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4949)
    
    wire \edb_top_inst/ceg_net24 , \edb_top_inst/la0/la_biu_inst/n1909 , 
        \edb_top_inst/la0/la_biu_inst/fifo_push , \edb_top_inst/n2823 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , \edb_top_inst/la0/la_biu_inst/fifo_rstn , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 , \edb_top_inst/~ceg_net27 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , \edb_top_inst/n2824 , 
        \edb_top_inst/n2825 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4581)
    
    wire \edb_top_inst/n2826 , \edb_top_inst/n2827 , \edb_top_inst/n2828 , 
        \edb_top_inst/n2829 , \edb_top_inst/n2830 , \edb_top_inst/n2831 , 
        \edb_top_inst/n2832 , \edb_top_inst/n2833 , \edb_top_inst/n2834 , 
        \edb_top_inst/n2835 , \edb_top_inst/n2836 , \edb_top_inst/n2837 , 
        \edb_top_inst/n2838 , \edb_top_inst/n2839 , \edb_top_inst/n2840 , 
        \edb_top_inst/n2841 , \edb_top_inst/n2842 , \edb_top_inst/n2843 , 
        \edb_top_inst/n2844 , \edb_top_inst/n2845 , \edb_top_inst/n2846 , 
        \edb_top_inst/n2847 , \edb_top_inst/n2848 , \edb_top_inst/n2849 , 
        \edb_top_inst/n2850 , \edb_top_inst/n2851 , \edb_top_inst/n2852 , 
        \edb_top_inst/n2853 , \edb_top_inst/n2854 , \edb_top_inst/n2855 , 
        \edb_top_inst/n2856 , \edb_top_inst/n2857 , \edb_top_inst/n2858 , 
        \edb_top_inst/n2859 , \edb_top_inst/n2860 , \edb_top_inst/n2861 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4581)
    
    wire \edb_top_inst/la0/n617 , \edb_top_inst/n2862 , \edb_top_inst/debug_hub_inst/n266 , 
        \edb_top_inst/debug_hub_inst/n95 , n2835;
    wire [7:0]rx_data;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(7)
    
    wire \uart_rx_inst/n925 , \uart_rx_inst/n896 , \uart_rx_inst/n899 , 
        ceg_net14, \uart_rx_inst/n924 , ceg_net32, \uart_rx_inst/n903 , 
        ceg_net26, \uart_rx_inst/n959 , \uart_rx_inst/n961 , \uart_rx_inst/n963 , 
        \uart_rx_inst/n965 , \uart_rx_inst/n967 , \uart_rx_inst/n969 , 
        \uart_rx_inst/n971 , \uart_rx_inst/n760 , \uart_rx_inst/n151 , 
        \uart_rx_inst/n955 , \uart_rx_inst/n767 , \uart_rx_inst/n770 , 
        \uart_rx_inst/n773 , \uart_rx_inst/n776 , \uart_rx_inst/n779 , 
        \uart_rx_inst/n782 , \uart_rx_inst/n785 , \uart_rx_inst/n788 , 
        \uart_rx_inst/n791 , \uart_rx_inst/n794 , \uart_rx_inst/n797 , 
        \uart_rx_inst/n800 , \uart_rx_inst/n803 , \uart_rx_inst/n806 , 
        \uart_rx_inst/n809 , \uart_rx_inst/n812 , \uart_rx_inst/n815 , 
        \uart_rx_inst/n818 , \uart_rx_inst/n821 , \uart_rx_inst/n824 , 
        \uart_rx_inst/n827 , \uart_rx_inst/n830 , \uart_rx_inst/n833 , 
        \uart_rx_inst/n836 , \uart_rx_inst/n839 , \uart_rx_inst/n842 , 
        \uart_rx_inst/n845 , \uart_rx_inst/n848 , \uart_rx_inst/n851 , 
        \uart_rx_inst/n854 , \uart_rx_inst/n857 , \uart_rx_inst/n861 , 
        \uart_rx_inst/n865 , \uart_tx_inst/n847 , \uart_tx_inst/n634 , 
        \uart_tx_inst/n851 , ceg_net28, \uart_tx_inst/n957 , \uart_tx_inst/n843 , 
        \uart_tx_inst/n716 , \uart_tx_inst/n719 , \uart_tx_inst/n722 , 
        \uart_tx_inst/n725 , \uart_tx_inst/n728 , \uart_tx_inst/n731 , 
        \uart_tx_inst/n734 , \uart_tx_inst/n737 , \uart_tx_inst/n810 , 
        \uart_tx_inst/n814 , \uart_tx_inst/n709 , \uart_tx_inst/LessThan_9/n18 , 
        \uart_tx_inst/n945 , \jtag_inst1_TCK~O , \clk~O , n2768, n2769, 
        n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
        n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
        n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
        n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
        n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
        n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
        n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, 
        n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
        n2834;
    
    EFX_LUT4 LUT__8043 (.I0(b[0]), .I1(a[0]), .O(n25)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(34)
    defparam LUT__8043.LUTMASK = 16'h6666;
    EFX_FF \b[0]~FF  (.D(rx_data[0]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \b[0]~FF .CLK_POLARITY = 1'b1;
    defparam \b[0]~FF .CE_POLARITY = 1'b1;
    defparam \b[0]~FF .SR_POLARITY = 1'b1;
    defparam \b[0]~FF .D_POLARITY = 1'b1;
    defparam \b[0]~FF .SR_SYNC = 1'b1;
    defparam \b[0]~FF .SR_VALUE = 1'b0;
    defparam \b[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \add_flag~FF  (.D(1'b1), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(add_flag)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \add_flag~FF .CLK_POLARITY = 1'b1;
    defparam \add_flag~FF .CE_POLARITY = 1'b1;
    defparam \add_flag~FF .SR_POLARITY = 1'b1;
    defparam \add_flag~FF .D_POLARITY = 1'b1;
    defparam \add_flag~FF .SR_SYNC = 1'b1;
    defparam \add_flag~FF .SR_VALUE = 1'b0;
    defparam \add_flag~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \send~FF  (.D(1'b1), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(send)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \send~FF .CLK_POLARITY = 1'b1;
    defparam \send~FF .CE_POLARITY = 1'b1;
    defparam \send~FF .SR_POLARITY = 1'b1;
    defparam \send~FF .D_POLARITY = 1'b1;
    defparam \send~FF .SR_SYNC = 1'b1;
    defparam \send~FF .SR_VALUE = 1'b0;
    defparam \send~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \sum[0]~FF  (.D(n25), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(sum[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \sum[0]~FF .CLK_POLARITY = 1'b1;
    defparam \sum[0]~FF .CE_POLARITY = 1'b1;
    defparam \sum[0]~FF .SR_POLARITY = 1'b1;
    defparam \sum[0]~FF .D_POLARITY = 1'b1;
    defparam \sum[0]~FF .SR_SYNC = 1'b1;
    defparam \sum[0]~FF .SR_VALUE = 1'b0;
    defparam \sum[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \carry~FF  (.D(n26[0]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(carry)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \carry~FF .CLK_POLARITY = 1'b1;
    defparam \carry~FF .CE_POLARITY = 1'b1;
    defparam \carry~FF .SR_POLARITY = 1'b1;
    defparam \carry~FF .D_POLARITY = 1'b1;
    defparam \carry~FF .SR_SYNC = 1'b1;
    defparam \carry~FF .SR_VALUE = 1'b0;
    defparam \carry~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[0]~FF  (.D(rx_data[4]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \a[0]~FF .CLK_POLARITY = 1'b1;
    defparam \a[0]~FF .CE_POLARITY = 1'b1;
    defparam \a[0]~FF .SR_POLARITY = 1'b1;
    defparam \a[0]~FF .D_POLARITY = 1'b1;
    defparam \a[0]~FF .SR_SYNC = 1'b1;
    defparam \a[0]~FF .SR_VALUE = 1'b0;
    defparam \a[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Data~FF  (.D(\uart_rx_inst/r_Rx_Data_R ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(102)
    defparam \uart_rx_inst/r_Rx_Data~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Data_R~FF  (.D(rx), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Data_R )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Data_R~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[0]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n925 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[0]~FF  (.D(\uart_rx_inst/n896 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/r_SM_Main [2]), .Q(\uart_rx_inst/r_SM_Main [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[0]~FF  (.D(\uart_rx_inst/n899 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_ready~FF  (.D(\uart_rx_inst/n924 ), .CE(ceg_net32), .CLK(\clk~O ), 
           .SR(1'b0), .Q(rx_ready)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \rx_ready~FF .CLK_POLARITY = 1'b1;
    defparam \rx_ready~FF .CE_POLARITY = 1'b0;
    defparam \rx_ready~FF .SR_POLARITY = 1'b1;
    defparam \rx_ready~FF .D_POLARITY = 1'b1;
    defparam \rx_ready~FF .SR_SYNC = 1'b1;
    defparam \rx_ready~FF .SR_VALUE = 1'b0;
    defparam \rx_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[0]~FF  (.D(\uart_rx_inst/n903 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[1]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n959 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[2]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n961 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[3]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n963 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[4]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n965 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[5]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n967 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[6]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n969 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[7]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n971 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[1]~FF  (.D(\uart_rx_inst/n760 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/r_SM_Main [2]), .Q(\uart_rx_inst/r_SM_Main [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[2]~FF  (.D(\uart_rx_inst/n151 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/n955 ), .Q(\uart_rx_inst/r_SM_Main [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[1]~FF  (.D(\uart_rx_inst/n767 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[2]~FF  (.D(\uart_rx_inst/n770 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[3]~FF  (.D(\uart_rx_inst/n773 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[4]~FF  (.D(\uart_rx_inst/n776 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[5]~FF  (.D(\uart_rx_inst/n779 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[6]~FF  (.D(\uart_rx_inst/n782 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[7]~FF  (.D(\uart_rx_inst/n785 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[8]~FF  (.D(\uart_rx_inst/n788 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[9]~FF  (.D(\uart_rx_inst/n791 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[10]~FF  (.D(\uart_rx_inst/n794 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[11]~FF  (.D(\uart_rx_inst/n797 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[12]~FF  (.D(\uart_rx_inst/n800 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[13]~FF  (.D(\uart_rx_inst/n803 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[14]~FF  (.D(\uart_rx_inst/n806 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[15]~FF  (.D(\uart_rx_inst/n809 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[16]~FF  (.D(\uart_rx_inst/n812 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[17]~FF  (.D(\uart_rx_inst/n815 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[18]~FF  (.D(\uart_rx_inst/n818 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[19]~FF  (.D(\uart_rx_inst/n821 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[20]~FF  (.D(\uart_rx_inst/n824 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[21]~FF  (.D(\uart_rx_inst/n827 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[22]~FF  (.D(\uart_rx_inst/n830 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[23]~FF  (.D(\uart_rx_inst/n833 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[24]~FF  (.D(\uart_rx_inst/n836 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[25]~FF  (.D(\uart_rx_inst/n839 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[26]~FF  (.D(\uart_rx_inst/n842 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[27]~FF  (.D(\uart_rx_inst/n845 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[28]~FF  (.D(\uart_rx_inst/n848 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[29]~FF  (.D(\uart_rx_inst/n851 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[30]~FF  (.D(\uart_rx_inst/n854 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[31]~FF  (.D(\uart_rx_inst/n857 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[1]~FF  (.D(\uart_rx_inst/n861 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[2]~FF  (.D(\uart_rx_inst/n865 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(176)
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[1]~FF  (.D(rx_data[1]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \b[1]~FF .CLK_POLARITY = 1'b1;
    defparam \b[1]~FF .CE_POLARITY = 1'b1;
    defparam \b[1]~FF .SR_POLARITY = 1'b1;
    defparam \b[1]~FF .D_POLARITY = 1'b1;
    defparam \b[1]~FF .SR_SYNC = 1'b1;
    defparam \b[1]~FF .SR_VALUE = 1'b0;
    defparam \b[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[2]~FF  (.D(rx_data[2]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \b[2]~FF .CLK_POLARITY = 1'b1;
    defparam \b[2]~FF .CE_POLARITY = 1'b1;
    defparam \b[2]~FF .SR_POLARITY = 1'b1;
    defparam \b[2]~FF .D_POLARITY = 1'b1;
    defparam \b[2]~FF .SR_SYNC = 1'b1;
    defparam \b[2]~FF .SR_VALUE = 1'b0;
    defparam \b[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[3]~FF  (.D(rx_data[3]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \b[3]~FF .CLK_POLARITY = 1'b1;
    defparam \b[3]~FF .CE_POLARITY = 1'b1;
    defparam \b[3]~FF .SR_POLARITY = 1'b1;
    defparam \b[3]~FF .D_POLARITY = 1'b1;
    defparam \b[3]~FF .SR_SYNC = 1'b1;
    defparam \b[3]~FF .SR_VALUE = 1'b0;
    defparam \b[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[0]~FF  (.D(\uart_tx_inst/n847 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_2~FF  (.D(\uart_tx_inst/n634 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(tx_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \tx_2~FF .CLK_POLARITY = 1'b1;
    defparam \tx_2~FF .CE_POLARITY = 1'b0;
    defparam \tx_2~FF .SR_POLARITY = 1'b1;
    defparam \tx_2~FF .D_POLARITY = 1'b0;
    defparam \tx_2~FF .SR_SYNC = 1'b1;
    defparam \tx_2~FF .SR_VALUE = 1'b0;
    defparam \tx_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[0]~FF  (.D(\uart_tx_inst/n851 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[0]~FF  (.D(sum[0]), .CE(\uart_tx_inst/n957 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[0]~FF  (.D(\uart_tx_inst/n843 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_tx_inst/r_SM_Main [2]), .Q(\uart_tx_inst/r_SM_Main [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[1]~FF  (.D(\uart_tx_inst/n716 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[2]~FF  (.D(\uart_tx_inst/n719 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[3]~FF  (.D(\uart_tx_inst/n722 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[4]~FF  (.D(\uart_tx_inst/n725 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[5]~FF  (.D(\uart_tx_inst/n728 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[6]~FF  (.D(\uart_tx_inst/n731 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[7]~FF  (.D(\uart_tx_inst/n734 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[8]~FF  (.D(\uart_tx_inst/n737 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[1]~FF  (.D(\uart_tx_inst/n810 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[2]~FF  (.D(\uart_tx_inst/n814 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[4]~FF  (.D(carry), .CE(\uart_tx_inst/n957 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[1]~FF  (.D(\uart_tx_inst/n709 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_tx_inst/r_SM_Main [2]), .Q(\uart_tx_inst/r_SM_Main [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[2]~FF  (.D(\uart_tx_inst/LessThan_9/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\uart_tx_inst/n945 ), .Q(\uart_tx_inst/r_SM_Main [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam \uart_tx_inst/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[1]~FF  (.D(rx_data[5]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \a[1]~FF .CLK_POLARITY = 1'b1;
    defparam \a[1]~FF .CE_POLARITY = 1'b1;
    defparam \a[1]~FF .SR_POLARITY = 1'b1;
    defparam \a[1]~FF .D_POLARITY = 1'b1;
    defparam \a[1]~FF .SR_SYNC = 1'b1;
    defparam \a[1]~FF .SR_VALUE = 1'b0;
    defparam \a[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[2]~FF  (.D(rx_data[6]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \a[2]~FF .CLK_POLARITY = 1'b1;
    defparam \a[2]~FF .CE_POLARITY = 1'b1;
    defparam \a[2]~FF .SR_POLARITY = 1'b1;
    defparam \a[2]~FF .D_POLARITY = 1'b1;
    defparam \a[2]~FF .SR_SYNC = 1'b1;
    defparam \a[2]~FF .SR_VALUE = 1'b0;
    defparam \a[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[3]~FF  (.D(rx_data[7]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(45)
    defparam \a[3]~FF .CLK_POLARITY = 1'b1;
    defparam \a[3]~FF .CE_POLARITY = 1'b1;
    defparam \a[3]~FF .SR_POLARITY = 1'b1;
    defparam \a[3]~FF .D_POLARITY = 1'b1;
    defparam \a[3]~FF .SR_SYNC = 1'b1;
    defparam \a[3]~FF .SR_VALUE = 1'b0;
    defparam \a[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1022 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1023 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1024 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1780 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [0]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3736)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n1998 [0]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [0]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2217 [0]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state [0]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3818)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/n2568 ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4128)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n2581 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n2568 ), .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4128)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(rx_ready), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n2581 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(rx_data[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3470 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3470 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(clk), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n4311 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(add_flag), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n5144 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n5144 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(rx), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n5977 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n6810 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n6810 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n6810 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(send), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n7643 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n7643 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n7643 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n8532 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n8532 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n8532 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n9429 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n9429 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n9429 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(a[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n10298 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n10298 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n10298 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n10313 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n10511 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF  (.D(b[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n11163 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n11163 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n11178 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n11376 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF  (.D(sum[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n12028 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n12028 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n12043 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n12241 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF  (.D(carry), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n12865 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n12865 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n12865 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF  (.D(tx_2), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n13698 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n13698 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr [64]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[8]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[9]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[10]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[11]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[12]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[13]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[14]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[15]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[16]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[17]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[18]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[19]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[20]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[21]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[22]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[23]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[24]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[25]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[26]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[27]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[28]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[29]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[30]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[31]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[32]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[33]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[34]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[35]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[36]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[37]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[38]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[39]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[40]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[41]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[42]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[43]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[44]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[45]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[46]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[47]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[48]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[49]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[50]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[51]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[52]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[53]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[54]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[55]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[56]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[57]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[58]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[59]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[60]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[61]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[62]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[63]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1595 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3679)
    defparam \edb_top_inst/la0/skip_count[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1728 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3692)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [1]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [2]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [3]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [4]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [5]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [6]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [7]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [8]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [9]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [10]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [11]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [12]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [13]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [14]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [15]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [16]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [17]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [18]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [19]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [20]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [21]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [22]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [23]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [24]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3726)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3736)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3736)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3736)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n1998 [1]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n1998 [2]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n1998 [3]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n1998 [4]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n1998 [5]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [1]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [2]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [3]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [4]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [5]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [6]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [7]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [8]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [9]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [10]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [11]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [12]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [13]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [14]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [15]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3763)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2217 [1]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2217 [2]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2217 [3]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2217 [4]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2217 [5]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2217 [6]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2217 [7]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2217 [8]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2217 [9]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2217 [10]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2217 [11]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2217 [12]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2217 [13]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2217 [14]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2217 [15]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2217 [16]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2217 [17]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2217 [18]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2217 [19]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2217 [20]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2217 [21]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2217 [22]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2217 [23]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2217 [24]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2217 [25]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2217 [26]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2217 [27]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2217 [28]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2217 [29]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2217 [30]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2217 [31]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2217 [32]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2217 [33]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2217 [34]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2217 [35]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2217 [36]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2217 [37]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2217 [38]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2217 [39]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2217 [40]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2217 [41]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2217 [42]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2217 [43]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2217 [44]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2217 [45]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2217 [46]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2217 [47]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2217 [48]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2217 [49]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2217 [50]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2217 [51]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2217 [52]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2217 [53]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2217 [54]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2217 [55]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2217 [56]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2217 [57]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2217 [58]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2217 [59]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2217 [60]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2217 [61]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2217 [62]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2217 [63]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3776)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state [1]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3818)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state [2]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3818)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state [3]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3818)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [0]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [1]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [2]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [3]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [4]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [5]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [6]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [7]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [8]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [9]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [10]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [11]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [12]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [13]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [14]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [15]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [16]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [17]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [18]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [19]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [20]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [21]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [22]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [23]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [24]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [25]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [26]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [27]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [28]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [29]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [30]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [31]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(288)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n2581 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF  (.D(rx_data[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF  (.D(rx_data[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF  (.D(rx_data[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF  (.D(rx_data[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF  (.D(rx_data[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF  (.D(rx_data[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF  (.D(rx_data[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3470 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n3485 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n3683 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n4311 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n4311 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n5144 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n5977 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n5977 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n8547 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n8745 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n9444 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n9642 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF  (.D(a[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF  (.D(a[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF  (.D(a[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n10313 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n10313 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n10313 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n10511 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n10511 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n10511 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF  (.D(b[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF  (.D(b[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF  (.D(b[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4155)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n7 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n11163 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n11178 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n11178 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n11178 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n11376 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n11376 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n11376 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/equal_9/n7 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n12028 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n12043 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n12043 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n12043 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n12241 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n12241 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n12241 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4279)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/equal_9/n7 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5676)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n13698 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5625)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5564)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n101 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5806)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[14]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[24]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[25]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[26]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[27]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[28]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[29]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[30]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[31]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[32]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [32]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[33]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [33]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[34]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [34]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[35]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [35]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[36]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [36]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[37]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [37]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[43]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4452)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [32]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [33]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [34]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [35]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [36]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [37]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [43]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4464)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [0]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/ts_trigger~FF  (.D(1'b1), .CE(\edb_top_inst/la0/trigger_skipper_n/n468 ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), .Q(\edb_top_inst/la0/ts_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/ts_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [1]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [2]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [3]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [4]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [5]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [6]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [7]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [8]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [9]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [10]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [11]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [12]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [13]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [14]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [15]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [16]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [17]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [18]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [19]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [20]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [21]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [22]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [23]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [24]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [25]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [26]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [27]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [28]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [29]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [30]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [31]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [32]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [33]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [34]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [35]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [36]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [37]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [38]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [39]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [40]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [41]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [42]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [43]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [44]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [45]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [46]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [47]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [48]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [49]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [50]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [51]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [52]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [53]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [54]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [55]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [56]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [57]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [58]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [59]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [60]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [61]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [62]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [63]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5881)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5292)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5092)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5092)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5092)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/ts_resetn~FF  (.D(\edb_top_inst/la0/la_biu_inst/n98 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/ts_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5092)
    defparam \edb_top_inst/la0/ts_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5313)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5328)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5328)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5328)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5338)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5351)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5351)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5351)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1319 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/n1902 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5475)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1284 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n19936 ), .Q(\edb_top_inst/la0/la_biu_inst/curr_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5292)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5292)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5292)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5092)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n370 ), 
           .CE(\edb_top_inst/ceg_net18 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5363)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter [15]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter [16]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter [17]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter [18]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter [19]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter [20]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter [21]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter [22]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter [23]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter [24]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n370 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5373)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [10]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [11]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [12]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [13]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [14]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [15]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [16]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [17]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [18]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [19]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [20]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [21]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [22]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [23]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [24]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [25]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [26]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [27]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [28]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [29]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [30]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [31]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [32]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [33]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [34]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[35]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [35]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[36]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [36]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[37]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [37]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[38]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [38]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[39]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [39]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[40]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [40]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[41]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [41]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [42]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[43]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [43]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[44]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [44]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1318 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5382)
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state [1]), 
           .CE(\edb_top_inst/ceg_net24 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5475)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt [0]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1909 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1909 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 [1]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [2]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [3]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [4]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [5]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [6]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [7]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [8]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [9]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [10]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4715)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [32]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [33]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [34]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [35]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [36]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [37]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [43]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4784)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [1]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [2]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [3]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [4]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [5]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [6]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [7]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [8]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [9]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [10]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr [65]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr [66]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr [67]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr [68]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr [69]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr [70]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr [71]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr [72]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr [73]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr [74]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr [75]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr [76]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3609)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n994 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(359)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(359)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(359)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(359)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr [64]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr [65]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr [66]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr [67]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr [68]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr [69]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr [70]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr [71]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr [72]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr [73]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr [74]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr [75]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr [76]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr [81]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(352)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \edb_top_inst/LUT__4339  (.I0(\edb_top_inst/la0/crc_data_out [24]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/la0/crc_data_out [31]), 
            .I3(\edb_top_inst/edb_user_dr [81]), .O(\edb_top_inst/n2056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4339 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4340  (.I0(\edb_top_inst/la0/crc_data_out [27]), 
            .I1(\edb_top_inst/edb_user_dr [77]), .I2(\edb_top_inst/la0/crc_data_out [28]), 
            .I3(\edb_top_inst/edb_user_dr [78]), .O(\edb_top_inst/n2057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4340 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4341  (.I0(\edb_top_inst/la0/crc_data_out [25]), 
            .I1(\edb_top_inst/edb_user_dr [75]), .I2(\edb_top_inst/la0/crc_data_out [26]), 
            .I3(\edb_top_inst/edb_user_dr [76]), .O(\edb_top_inst/n2058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4341 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4342  (.I0(\edb_top_inst/n2055 ), .I1(\edb_top_inst/n2056 ), 
            .I2(\edb_top_inst/n2057 ), .I3(\edb_top_inst/n2058 ), .O(\edb_top_inst/n2059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4342 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4343  (.I0(\edb_top_inst/la0/crc_data_out [16]), 
            .I1(\edb_top_inst/edb_user_dr [66]), .I2(\edb_top_inst/la0/crc_data_out [23]), 
            .I3(\edb_top_inst/edb_user_dr [73]), .O(\edb_top_inst/n2060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4343 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4344  (.I0(\edb_top_inst/la0/crc_data_out [19]), 
            .I1(\edb_top_inst/edb_user_dr [69]), .I2(\edb_top_inst/la0/crc_data_out [20]), 
            .I3(\edb_top_inst/edb_user_dr [70]), .O(\edb_top_inst/n2061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4344 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4345  (.I0(\edb_top_inst/la0/crc_data_out [17]), 
            .I1(\edb_top_inst/edb_user_dr [67]), .I2(\edb_top_inst/la0/crc_data_out [18]), 
            .I3(\edb_top_inst/edb_user_dr [68]), .O(\edb_top_inst/n2062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4345 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4346  (.I0(\edb_top_inst/la0/crc_data_out [21]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/la0/crc_data_out [22]), 
            .I3(\edb_top_inst/edb_user_dr [72]), .O(\edb_top_inst/n2063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4346 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4347  (.I0(\edb_top_inst/n2060 ), .I1(\edb_top_inst/n2061 ), 
            .I2(\edb_top_inst/n2062 ), .I3(\edb_top_inst/n2063 ), .O(\edb_top_inst/n2064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4347 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4348  (.I0(\edb_top_inst/la0/crc_data_out [10]), 
            .I1(\edb_top_inst/edb_user_dr [60]), .I2(\edb_top_inst/la0/crc_data_out [11]), 
            .I3(\edb_top_inst/edb_user_dr [61]), .O(\edb_top_inst/n2065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4348 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4349  (.I0(\edb_top_inst/la0/crc_data_out [8]), 
            .I1(\edb_top_inst/edb_user_dr [58]), .I2(\edb_top_inst/la0/crc_data_out [9]), 
            .I3(\edb_top_inst/edb_user_dr [59]), .O(\edb_top_inst/n2066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4349 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4350  (.I0(\edb_top_inst/la0/crc_data_out [12]), 
            .I1(\edb_top_inst/edb_user_dr [62]), .I2(\edb_top_inst/la0/crc_data_out [13]), 
            .I3(\edb_top_inst/edb_user_dr [63]), .O(\edb_top_inst/n2067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4350 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4351  (.I0(\edb_top_inst/la0/crc_data_out [7]), 
            .I1(\edb_top_inst/edb_user_dr [57]), .I2(\edb_top_inst/la0/crc_data_out [14]), 
            .I3(\edb_top_inst/edb_user_dr [64]), .O(\edb_top_inst/n2068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4351 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4352  (.I0(\edb_top_inst/n2065 ), .I1(\edb_top_inst/n2066 ), 
            .I2(\edb_top_inst/n2067 ), .I3(\edb_top_inst/n2068 ), .O(\edb_top_inst/n2069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4352 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4353  (.I0(\edb_top_inst/la0/crc_data_out [2]), 
            .I1(\edb_top_inst/edb_user_dr [52]), .I2(\edb_top_inst/la0/crc_data_out [3]), 
            .I3(\edb_top_inst/edb_user_dr [53]), .O(\edb_top_inst/n2070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4353 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4354  (.I0(\edb_top_inst/la0/crc_data_out [4]), 
            .I1(\edb_top_inst/edb_user_dr [54]), .I2(\edb_top_inst/la0/crc_data_out [5]), 
            .I3(\edb_top_inst/edb_user_dr [55]), .O(\edb_top_inst/n2071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4354 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4355  (.I0(\edb_top_inst/la0/crc_data_out [6]), 
            .I1(\edb_top_inst/edb_user_dr [56]), .I2(\edb_top_inst/la0/crc_data_out [15]), 
            .I3(\edb_top_inst/edb_user_dr [65]), .O(\edb_top_inst/n2072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4355 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4356  (.I0(\edb_top_inst/la0/crc_data_out [0]), 
            .I1(\edb_top_inst/edb_user_dr [50]), .I2(\edb_top_inst/la0/crc_data_out [1]), 
            .I3(\edb_top_inst/edb_user_dr [51]), .O(\edb_top_inst/n2073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4356 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4357  (.I0(\edb_top_inst/n2070 ), .I1(\edb_top_inst/n2071 ), 
            .I2(\edb_top_inst/n2072 ), .I3(\edb_top_inst/n2073 ), .O(\edb_top_inst/n2074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4357 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4358  (.I0(\edb_top_inst/n2059 ), .I1(\edb_top_inst/n2064 ), 
            .I2(\edb_top_inst/n2069 ), .I3(\edb_top_inst/n2074 ), .O(\edb_top_inst/n2075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4358 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4359  (.I0(\edb_top_inst/la0/bit_count [3]), 
            .I1(\edb_top_inst/la0/bit_count [4]), .I2(\edb_top_inst/la0/bit_count [5]), 
            .I3(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n2076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4359 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4360  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/la0/bit_count [1]), .I2(\edb_top_inst/la0/bit_count [2]), 
            .I3(\edb_top_inst/n2076 ), .O(\edb_top_inst/n2077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4360 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4361  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n2077 ), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n2078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4361 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4362  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/la0/module_state [0]), .O(\edb_top_inst/n2079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4362 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4363  (.I0(\edb_top_inst/n2078 ), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(\edb_top_inst/n2079 ), .I3(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n2080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4363 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4364  (.I0(\edb_top_inst/n2075 ), .I1(\edb_top_inst/la0/crc_data_out [0]), 
            .I2(\edb_top_inst/n2080 ), .O(\edb_top_inst/n2081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4364 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4365  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg [0]), .I2(\edb_top_inst/n2080 ), 
            .O(\edb_top_inst/n2082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4365 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4366  (.I0(\edb_top_inst/la0/word_count [0]), 
            .I1(\edb_top_inst/la0/word_count [1]), .I2(\edb_top_inst/la0/word_count [2]), 
            .I3(\edb_top_inst/la0/word_count [3]), .O(\edb_top_inst/n2083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4366 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4367  (.I0(\edb_top_inst/la0/word_count [4]), 
            .I1(\edb_top_inst/la0/word_count [5]), .I2(\edb_top_inst/la0/word_count [6]), 
            .I3(\edb_top_inst/la0/word_count [7]), .O(\edb_top_inst/n2084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4367 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4368  (.I0(\edb_top_inst/la0/word_count [12]), 
            .I1(\edb_top_inst/la0/word_count [13]), .I2(\edb_top_inst/la0/word_count [14]), 
            .I3(\edb_top_inst/la0/word_count [15]), .O(\edb_top_inst/n2085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4368 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4369  (.I0(\edb_top_inst/la0/word_count [8]), 
            .I1(\edb_top_inst/la0/word_count [9]), .I2(\edb_top_inst/la0/word_count [10]), 
            .I3(\edb_top_inst/la0/word_count [11]), .O(\edb_top_inst/n2086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4369 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4370  (.I0(\edb_top_inst/n2083 ), .I1(\edb_top_inst/n2084 ), 
            .I2(\edb_top_inst/n2085 ), .I3(\edb_top_inst/n2086 ), .O(\edb_top_inst/n2087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4370 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4371  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n2088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4371 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4372  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n2087 ), 
            .I2(\edb_top_inst/n2088 ), .O(\edb_top_inst/n2089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4372 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4373  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [3]), .O(\edb_top_inst/la0/n619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4373 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4374  (.I0(\edb_top_inst/la0/opcode [3]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [0]), .O(\edb_top_inst/la0/n618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4374 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4375  (.I0(\edb_top_inst/la0/n619 ), .I1(\edb_top_inst/la0/n618 ), 
            .I2(\edb_top_inst/la0/bit_count [5]), .I3(\edb_top_inst/la0/bit_count [4]), 
            .O(\edb_top_inst/n2090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4375 .LUTMASK = 16'h53fe;
    EFX_LUT4 \edb_top_inst/LUT__4376  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [3]), .O(\edb_top_inst/n2091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4376 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4377  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/la0/bit_count [1]), .I2(\edb_top_inst/la0/bit_count [2]), 
            .I3(\edb_top_inst/n2091 ), .O(\edb_top_inst/n2092 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4377 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__4378  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [3]), .O(\edb_top_inst/n2093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4378 .LUTMASK = 16'hfe3f;
    EFX_LUT4 \edb_top_inst/LUT__4379  (.I0(\edb_top_inst/n2090 ), .I1(\edb_top_inst/n2092 ), 
            .I2(\edb_top_inst/la0/bit_count [3]), .I3(\edb_top_inst/n2093 ), 
            .O(\edb_top_inst/n2094 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4379 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__4380  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .I2(\edb_top_inst/n2094 ), 
            .O(\edb_top_inst/n2095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4380 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__4381  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n2096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4381 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4382  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n2097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4382 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4383  (.I0(\edb_top_inst/n2096 ), .I1(\edb_top_inst/n2087 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n2097 ), .O(\edb_top_inst/n2098 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4383 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4384  (.I0(\edb_top_inst/n2095 ), .I1(\edb_top_inst/n2089 ), 
            .I2(\edb_top_inst/n2098 ), .O(\edb_top_inst/la0/module_next_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4384 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4385  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n2099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4385 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4386  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg [1]), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg [2]), .I2(\edb_top_inst/debug_hub_inst/module_id_reg [3]), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg [0]), .O(\edb_top_inst/n2100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4386 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4387  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n2100 ), 
            .O(\edb_top_inst/n2101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4387 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4388  (.I0(\edb_top_inst/n2087 ), .I1(\edb_top_inst/n2101 ), 
            .I2(\edb_top_inst/la0/module_state [0]), .I3(\edb_top_inst/la0/module_state [1]), 
            .O(\edb_top_inst/n2102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4388 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4389  (.I0(\edb_top_inst/n2087 ), .I1(\edb_top_inst/n2099 ), 
            .I2(\edb_top_inst/n2094 ), .I3(\edb_top_inst/n2102 ), .O(\edb_top_inst/n2103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4389 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4390  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n2104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4390 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4391  (.I0(\edb_top_inst/n2099 ), .I1(\edb_top_inst/edb_user_dr [81]), 
            .I2(\edb_top_inst/n2100 ), .I3(\edb_top_inst/la0/module_state [1]), 
            .O(\edb_top_inst/n2105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4391 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4392  (.I0(\edb_top_inst/n2094 ), .I1(\edb_top_inst/n2087 ), 
            .I2(\edb_top_inst/n2104 ), .I3(\edb_top_inst/n2105 ), .O(\edb_top_inst/n2106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4392 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4393  (.I0(\edb_top_inst/n2087 ), .I1(\edb_top_inst/la0/module_state [1]), 
            .I2(\edb_top_inst/la0/module_state [0]), .I3(\edb_top_inst/n2077 ), 
            .O(\edb_top_inst/n2107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4393 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4394  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n2108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4394 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4395  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n2109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4395 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4396  (.I0(\edb_top_inst/n2100 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n2109 ), .I3(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n2110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4396 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__4397  (.I0(\edb_top_inst/edb_user_dr [77]), 
            .I1(\edb_top_inst/edb_user_dr [78]), .I2(\edb_top_inst/edb_user_dr [79]), 
            .I3(\edb_top_inst/edb_user_dr [80]), .O(\edb_top_inst/n2111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4397 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4398  (.I0(\edb_top_inst/edb_user_dr [81]), 
            .I1(jtag_inst1_UPDATE), .O(\edb_top_inst/n2112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4398 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4399  (.I0(\edb_top_inst/n2111 ), .I1(\edb_top_inst/n2100 ), 
            .I2(\edb_top_inst/n2112 ), .I3(\edb_top_inst/n2096 ), .O(\edb_top_inst/n2113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4399 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4400  (.I0(\edb_top_inst/n2110 ), .I1(\edb_top_inst/la0/module_state [1]), 
            .I2(\edb_top_inst/n2113 ), .I3(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n2114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4400 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__4401  (.I0(\edb_top_inst/n2107 ), .I1(\edb_top_inst/n2108 ), 
            .I2(\edb_top_inst/n2114 ), .I3(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n2115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4401 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__4402  (.I0(\edb_top_inst/n2106 ), .I1(\edb_top_inst/n2103 ), 
            .I2(\edb_top_inst/n2088 ), .I3(\edb_top_inst/n2115 ), .O(\edb_top_inst/la0/module_next_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4402 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__4403  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/la0/module_next_state [3]), .I2(\edb_top_inst/la0/module_state [0]), 
            .I3(\edb_top_inst/n2097 ), .O(\edb_top_inst/n2116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4403 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4404  (.I0(\edb_top_inst/n2082 ), .I1(\edb_top_inst/n2081 ), 
            .I2(\edb_top_inst/n2116 ), .I3(\edb_top_inst/n2100 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4404 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4405  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [40]), .O(\edb_top_inst/la0/n1022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4405 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4406  (.I0(\edb_top_inst/edb_user_dr [75]), 
            .I1(\edb_top_inst/edb_user_dr [76]), .O(\edb_top_inst/n2117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4406 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4407  (.I0(\edb_top_inst/edb_user_dr [73]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/n2117 ), 
            .O(\edb_top_inst/n2118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4407 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4408  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/edb_user_dr [72]), 
            .O(\edb_top_inst/n2119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4408 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4409  (.I0(\edb_top_inst/n2118 ), .I1(\edb_top_inst/n2119 ), 
            .O(\edb_top_inst/n2120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4409 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4410  (.I0(\edb_top_inst/edb_user_dr [78]), 
            .I1(\edb_top_inst/edb_user_dr [77]), .I2(\edb_top_inst/edb_user_dr [80]), 
            .O(\edb_top_inst/n2121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4410 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4411  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .I2(\edb_top_inst/la0/module_state [2]), 
            .I3(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n2122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4411 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4412  (.I0(\edb_top_inst/n2100 ), .I1(\edb_top_inst/n2112 ), 
            .I2(\edb_top_inst/n2121 ), .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4412 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4413  (.I0(\edb_top_inst/edb_user_dr [68]), 
            .I1(\edb_top_inst/edb_user_dr [69]), .I2(\edb_top_inst/edb_user_dr [79]), 
            .I3(\edb_top_inst/la0/regsel_ld_en ), .O(\edb_top_inst/n2123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4413 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4414  (.I0(\edb_top_inst/edb_user_dr [66]), 
            .I1(\edb_top_inst/edb_user_dr [67]), .I2(\edb_top_inst/n2123 ), 
            .O(\edb_top_inst/n2124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4414 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4415  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n2124 ), 
            .O(\edb_top_inst/n2125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4415 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4416  (.I0(\edb_top_inst/n2120 ), .I1(\edb_top_inst/n2125 ), 
            .O(\edb_top_inst/la0/n994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4416 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4417  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/la0/n994 ), .O(\edb_top_inst/ceg_net2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4417 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4418  (.I0(\edb_top_inst/edb_user_dr [65]), 
            .I1(\edb_top_inst/edb_user_dr [64]), .I2(\edb_top_inst/n2124 ), 
            .O(\edb_top_inst/n2126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4418 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4419  (.I0(\edb_top_inst/n2120 ), .I1(\edb_top_inst/n2126 ), 
            .O(\edb_top_inst/la0/n1078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4419 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4420  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [41]), .O(\edb_top_inst/la0/n1023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4420 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4421  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [42]), .O(\edb_top_inst/la0/n1024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4421 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4422  (.I0(\edb_top_inst/n2120 ), .I1(\edb_top_inst/n2123 ), 
            .O(\edb_top_inst/n2127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4422 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4423  (.I0(\edb_top_inst/edb_user_dr [66]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n2127 ), 
            .O(\edb_top_inst/n2128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4423 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4424  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [67]), .I2(\edb_top_inst/n2128 ), 
            .O(\edb_top_inst/la0/n1595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4424 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4425  (.I0(\edb_top_inst/edb_user_dr [67]), 
            .I1(\edb_top_inst/edb_user_dr [64]), .I2(\edb_top_inst/n2128 ), 
            .O(\edb_top_inst/la0/n1728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4425 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4426  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/edb_user_dr [67]), 
            .I3(\edb_top_inst/edb_user_dr [66]), .O(\edb_top_inst/n2129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4426 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4427  (.I0(\edb_top_inst/edb_user_dr [63]), 
            .I1(\edb_top_inst/n2127 ), .I2(\edb_top_inst/n2129 ), .O(\edb_top_inst/la0/n1780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4427 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4428  (.I0(\edb_top_inst/la0/address_counter [0]), 
            .I1(\edb_top_inst/la0/address_counter [1]), .I2(\edb_top_inst/la0/address_counter [2]), 
            .I3(\edb_top_inst/la0/address_counter [6]), .O(\edb_top_inst/n2130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4428 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4429  (.I0(\edb_top_inst/la0/address_counter [3]), 
            .I1(\edb_top_inst/la0/address_counter [4]), .I2(\edb_top_inst/la0/address_counter [5]), 
            .I3(\edb_top_inst/la0/address_counter [14]), .O(\edb_top_inst/n2131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4429 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4430  (.I0(\edb_top_inst/la0/address_counter [7]), 
            .I1(\edb_top_inst/la0/address_counter [8]), .I2(\edb_top_inst/la0/address_counter [9]), 
            .I3(\edb_top_inst/la0/address_counter [10]), .O(\edb_top_inst/n2132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4430 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4431  (.I0(\edb_top_inst/la0/address_counter [11]), 
            .I1(\edb_top_inst/la0/address_counter [12]), .I2(\edb_top_inst/la0/address_counter [13]), 
            .O(\edb_top_inst/n2133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4431 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4432  (.I0(\edb_top_inst/n2130 ), .I1(\edb_top_inst/n2131 ), 
            .I2(\edb_top_inst/n2132 ), .I3(\edb_top_inst/n2133 ), .O(\edb_top_inst/n2134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4432 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4433  (.I0(\edb_top_inst/n2134 ), .I1(\edb_top_inst/la0/n1837 [0]), 
            .I2(\edb_top_inst/edb_user_dr [45]), .I3(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4433 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4434  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/n2087 ), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/la0/module_state [0]), .O(\edb_top_inst/n2135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4434 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__4435  (.I0(\edb_top_inst/la0/word_count [8]), 
            .I1(\edb_top_inst/la0/word_count [9]), .I2(\edb_top_inst/la0/word_count [10]), 
            .O(\edb_top_inst/n2136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4435 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4436  (.I0(\edb_top_inst/la0/word_count [11]), 
            .I1(\edb_top_inst/n2084 ), .I2(\edb_top_inst/n2136 ), .I3(\edb_top_inst/n2085 ), 
            .O(\edb_top_inst/n2137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4436 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4437  (.I0(\edb_top_inst/la0/word_count [1]), 
            .I1(\edb_top_inst/la0/word_count [2]), .I2(\edb_top_inst/la0/word_count [3]), 
            .I3(\edb_top_inst/n2137 ), .O(\edb_top_inst/n2138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4437 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4438  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [2]), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n2139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4438 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4439  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(\edb_top_inst/n2139 ), 
            .O(\edb_top_inst/n2140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4439 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4440  (.I0(\edb_top_inst/n2140 ), .I1(\edb_top_inst/n2138 ), 
            .I2(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n2141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4440 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4441  (.I0(\edb_top_inst/n2138 ), .I1(\edb_top_inst/la0/module_state [1]), 
            .I2(\edb_top_inst/la0/module_state [0]), .I3(\edb_top_inst/n2094 ), 
            .O(\edb_top_inst/n2142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4441 .LUTMASK = 16'hc100;
    EFX_LUT4 \edb_top_inst/LUT__4442  (.I0(\edb_top_inst/n2142 ), .I1(\edb_top_inst/la0/module_state [2]), 
            .I2(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n2143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4442 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4443  (.I0(\edb_top_inst/n2097 ), .I1(\edb_top_inst/n2096 ), 
            .O(\edb_top_inst/n2144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4443 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4444  (.I0(\edb_top_inst/n2135 ), .I1(\edb_top_inst/n2141 ), 
            .I2(\edb_top_inst/n2143 ), .I3(\edb_top_inst/n2144 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4444 .LUTMASK = 16'hffb0;
    EFX_LUT4 \edb_top_inst/LUT__4445  (.I0(\edb_top_inst/la0/opcode [1]), 
            .I1(\edb_top_inst/la0/opcode [3]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [0]), .O(\edb_top_inst/la0/n616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4445 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4446  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4446 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4447  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/n2096 ), .O(\edb_top_inst/n2145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4447 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4448  (.I0(\edb_top_inst/n2095 ), .I1(\edb_top_inst/la0/module_state [2]), 
            .I2(\edb_top_inst/n2140 ), .O(\edb_top_inst/n2146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4448 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4449  (.I0(\edb_top_inst/n2146 ), .I1(\edb_top_inst/la0/module_next_state [0]), 
            .I2(\edb_top_inst/n2145 ), .I3(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n2147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0d5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4449 .LUTMASK = 16'hf0d5;
    EFX_LUT4 \edb_top_inst/LUT__4450  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/n2147 ), .O(\edb_top_inst/la0/n1998 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4450 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4451  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [2]), .I2(\edb_top_inst/la0/module_state [3]), 
            .I3(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n2148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4451 .LUTMASK = 16'h1800;
    EFX_LUT4 \edb_top_inst/LUT__4452  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/n2088 ), .O(\edb_top_inst/n2149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4452 .LUTMASK = 16'he300;
    EFX_LUT4 \edb_top_inst/LUT__4453  (.I0(\edb_top_inst/n2148 ), .I1(\edb_top_inst/n2149 ), 
            .I2(\edb_top_inst/n2147 ), .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4453 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4454  (.I0(\edb_top_inst/edb_user_dr [29]), 
            .I1(\edb_top_inst/la0/word_count [0]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_word_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4454 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4455  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/la0/module_state [1]), .I2(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n2150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4455 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4456  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/n2150 ), .I2(\edb_top_inst/n2094 ), .I3(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n2151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf15, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4456 .LUTMASK = 16'hcf15;
    EFX_LUT4 \edb_top_inst/LUT__4457  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/n2151 ), 
            .I2(\edb_top_inst/n2088 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4457 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4458  (.I0(\edb_top_inst/la0/internal_register_select [9]), 
            .I1(\edb_top_inst/la0/internal_register_select [10]), .I2(\edb_top_inst/la0/internal_register_select [11]), 
            .I3(\edb_top_inst/la0/internal_register_select [12]), .O(\edb_top_inst/n2152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4458 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4459  (.I0(\edb_top_inst/la0/internal_register_select [2]), 
            .I1(\edb_top_inst/la0/internal_register_select [6]), .I2(\edb_top_inst/la0/internal_register_select [7]), 
            .I3(\edb_top_inst/la0/internal_register_select [8]), .O(\edb_top_inst/n2153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4459 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4460  (.I0(\edb_top_inst/la0/internal_register_select [4]), 
            .I1(\edb_top_inst/la0/internal_register_select [5]), .O(\edb_top_inst/n2154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4460 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4461  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/la0/internal_register_select [1]), .I2(\edb_top_inst/la0/internal_register_select [3]), 
            .O(\edb_top_inst/n2155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4461 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4462  (.I0(\edb_top_inst/n2152 ), .I1(\edb_top_inst/n2153 ), 
            .I2(\edb_top_inst/n2154 ), .I3(\edb_top_inst/n2155 ), .O(\edb_top_inst/n2156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4462 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4463  (.I0(\edb_top_inst/la0/la_trig_mask [0]), 
            .I1(\edb_top_inst/la0/internal_register_select [0]), .O(\edb_top_inst/n2157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4463 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4464  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/la0/internal_register_select [4]), .I2(\edb_top_inst/la0/internal_register_select [5]), 
            .O(\edb_top_inst/n2158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4464 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4465  (.I0(\edb_top_inst/la0/internal_register_select [1]), 
            .I1(\edb_top_inst/n2152 ), .I2(\edb_top_inst/n2153 ), .I3(\edb_top_inst/n2158 ), 
            .O(\edb_top_inst/n2159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4465 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4466  (.I0(\edb_top_inst/n2157 ), .I1(\edb_top_inst/n2159 ), 
            .I2(\edb_top_inst/la0/skip_count [0]), .I3(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4466 .LUTMASK = 16'h0bbb;
    EFX_LUT4 \edb_top_inst/LUT__4467  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4467 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4468  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/n2162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h13f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4468 .LUTMASK = 16'h13f8;
    EFX_LUT4 \edb_top_inst/LUT__4469  (.I0(\edb_top_inst/n2162 ), .I1(\edb_top_inst/n2161 ), 
            .O(\edb_top_inst/n2163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4469 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4470  (.I0(\edb_top_inst/n2096 ), .I1(\edb_top_inst/n2094 ), 
            .I2(\edb_top_inst/n2088 ), .I3(\edb_top_inst/n2140 ), .O(\edb_top_inst/n2164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4470 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__4471  (.I0(\edb_top_inst/n2163 ), .I1(\edb_top_inst/n2160 ), 
            .I2(\edb_top_inst/la0/data_from_biu [0]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4471 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4472  (.I0(\edb_top_inst/n2096 ), .I1(\edb_top_inst/n2101 ), 
            .I2(\edb_top_inst/n2140 ), .O(\edb_top_inst/n2166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4472 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4473  (.I0(\edb_top_inst/n2096 ), .I1(\edb_top_inst/n2094 ), 
            .I2(\edb_top_inst/n2166 ), .I3(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n2167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4473 .LUTMASK = 16'h77f0;
    EFX_LUT4 \edb_top_inst/LUT__4474  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/n2167 ), .O(\edb_top_inst/n2168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4474 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4475  (.I0(\edb_top_inst/n2165 ), .I1(\edb_top_inst/la0/data_out_shift_reg [1]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4475 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4476  (.I0(\edb_top_inst/n2100 ), .I1(jtag_inst1_SHIFT), 
            .I2(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n2169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4476 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4477  (.I0(\edb_top_inst/n2169 ), .I1(\edb_top_inst/n2096 ), 
            .I2(\edb_top_inst/n2167 ), .I3(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/ceg_net8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4477 .LUTMASK = 16'hffb0;
    EFX_LUT4 \edb_top_inst/LUT__4478  (.I0(jtag_inst1_RESET), .I1(\edb_top_inst/la0/la_soft_reset_in ), 
            .O(\edb_top_inst/la0/n2568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4478 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4479  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [72]), .I2(\edb_top_inst/edb_user_dr [71]), 
            .O(\edb_top_inst/n2170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4479 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4480  (.I0(\edb_top_inst/n2118 ), .I1(\edb_top_inst/n2125 ), 
            .O(\edb_top_inst/n2171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4480 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4481  (.I0(\edb_top_inst/n2170 ), .I1(\edb_top_inst/n2171 ), 
            .O(\edb_top_inst/la0/n2581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4481 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4482  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/edb_user_dr [72]), 
            .O(\edb_top_inst/n2172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4482 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4483  (.I0(\edb_top_inst/n2118 ), .I1(\edb_top_inst/n2172 ), 
            .O(\edb_top_inst/n2173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4483 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4484  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2173 ), 
            .O(\edb_top_inst/la0/n3470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4484 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4485  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2173 ), 
            .O(\edb_top_inst/la0/n3485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4485 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4486  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n2124 ), 
            .O(\edb_top_inst/n2174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4486 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4487  (.I0(\edb_top_inst/n2173 ), .I1(\edb_top_inst/n2174 ), 
            .O(\edb_top_inst/la0/n3683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4487 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4488  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/edb_user_dr [72]), 
            .I3(\edb_top_inst/n2171 ), .O(\edb_top_inst/la0/n4311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4488 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4489  (.I0(\edb_top_inst/edb_user_dr [74]), 
            .I1(\edb_top_inst/edb_user_dr [73]), .I2(\edb_top_inst/n2117 ), 
            .I3(\edb_top_inst/n2125 ), .O(\edb_top_inst/n2175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4489 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4490  (.I0(\edb_top_inst/n2119 ), .I1(\edb_top_inst/n2175 ), 
            .O(\edb_top_inst/la0/n5144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4490 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4491  (.I0(\edb_top_inst/n2170 ), .I1(\edb_top_inst/n2175 ), 
            .O(\edb_top_inst/la0/n5977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4491 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4492  (.I0(\edb_top_inst/n2172 ), .I1(\edb_top_inst/n2175 ), 
            .O(\edb_top_inst/la0/n6810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4492 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4493  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/edb_user_dr [72]), 
            .I3(\edb_top_inst/n2175 ), .O(\edb_top_inst/la0/n7643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4493 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4494  (.I0(\edb_top_inst/edb_user_dr [73]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/n2117 ), 
            .O(\edb_top_inst/n2176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4494 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4495  (.I0(\edb_top_inst/n2119 ), .I1(\edb_top_inst/n2176 ), 
            .O(\edb_top_inst/n2177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4495 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4496  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2177 ), 
            .O(\edb_top_inst/la0/n8532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4496 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4497  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2177 ), 
            .O(\edb_top_inst/la0/n8547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4497 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4498  (.I0(\edb_top_inst/n2174 ), .I1(\edb_top_inst/n2177 ), 
            .O(\edb_top_inst/la0/n8745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4498 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4499  (.I0(\edb_top_inst/n2170 ), .I1(\edb_top_inst/n2176 ), 
            .O(\edb_top_inst/n2178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4499 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4500  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2178 ), 
            .O(\edb_top_inst/la0/n9429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4500 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4501  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2178 ), 
            .O(\edb_top_inst/la0/n9444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4501 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4502  (.I0(\edb_top_inst/n2174 ), .I1(\edb_top_inst/n2178 ), 
            .O(\edb_top_inst/la0/n9642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4502 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4503  (.I0(\edb_top_inst/n2172 ), .I1(\edb_top_inst/n2176 ), 
            .O(\edb_top_inst/n2179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4503 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4504  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2179 ), 
            .O(\edb_top_inst/la0/n10298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4504 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4505  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2179 ), 
            .O(\edb_top_inst/la0/n10313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4505 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4506  (.I0(\edb_top_inst/n2174 ), .I1(\edb_top_inst/n2179 ), 
            .O(\edb_top_inst/la0/n10511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4506 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4507  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/edb_user_dr [72]), 
            .I3(\edb_top_inst/n2176 ), .O(\edb_top_inst/n2180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4507 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4508  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2180 ), 
            .O(\edb_top_inst/la0/n11163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4508 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4509  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2180 ), 
            .O(\edb_top_inst/la0/n11178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4509 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4510  (.I0(\edb_top_inst/n2174 ), .I1(\edb_top_inst/n2180 ), 
            .O(\edb_top_inst/la0/n11376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4510 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4511  (.I0(\edb_top_inst/edb_user_dr [73]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/n2117 ), 
            .I3(\edb_top_inst/n2119 ), .O(\edb_top_inst/n2181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4511 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4512  (.I0(\edb_top_inst/n2125 ), .I1(\edb_top_inst/n2181 ), 
            .O(\edb_top_inst/la0/n12028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4512 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4513  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2181 ), 
            .O(\edb_top_inst/la0/n12043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4513 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4514  (.I0(\edb_top_inst/n2174 ), .I1(\edb_top_inst/n2181 ), 
            .O(\edb_top_inst/la0/n12241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4514 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4515  (.I0(\edb_top_inst/edb_user_dr [73]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/n2117 ), 
            .I3(\edb_top_inst/n2125 ), .O(\edb_top_inst/n2182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4515 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4516  (.I0(\edb_top_inst/n2170 ), .I1(\edb_top_inst/n2182 ), 
            .O(\edb_top_inst/la0/n12865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4516 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4517  (.I0(\edb_top_inst/n2172 ), .I1(\edb_top_inst/n2182 ), 
            .O(\edb_top_inst/la0/n13698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4517 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4518  (.I0(\edb_top_inst/n2134 ), .I1(\edb_top_inst/la0/n1837 [1]), 
            .I2(\edb_top_inst/edb_user_dr [46]), .I3(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4518 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4519  (.I0(\edb_top_inst/n2134 ), .I1(\edb_top_inst/la0/n1837 [2]), 
            .I2(\edb_top_inst/edb_user_dr [47]), .I3(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4519 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4520  (.I0(\edb_top_inst/n2134 ), .I1(\edb_top_inst/la0/n1837 [3]), 
            .I2(\edb_top_inst/edb_user_dr [48]), .I3(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4520 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4521  (.I0(\edb_top_inst/edb_user_dr [49]), 
            .I1(\edb_top_inst/la0/n1837 [4]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4521 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4522  (.I0(\edb_top_inst/edb_user_dr [50]), 
            .I1(\edb_top_inst/la0/n1837 [5]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4522 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4523  (.I0(\edb_top_inst/edb_user_dr [51]), 
            .I1(\edb_top_inst/la0/n1837 [6]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4523 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4524  (.I0(\edb_top_inst/edb_user_dr [52]), 
            .I1(\edb_top_inst/la0/n1837 [7]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4524 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4525  (.I0(\edb_top_inst/edb_user_dr [53]), 
            .I1(\edb_top_inst/la0/n1837 [8]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4525 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4526  (.I0(\edb_top_inst/edb_user_dr [54]), 
            .I1(\edb_top_inst/la0/n1837 [9]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4526 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4527  (.I0(\edb_top_inst/edb_user_dr [55]), 
            .I1(\edb_top_inst/la0/n1837 [10]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4527 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4528  (.I0(\edb_top_inst/edb_user_dr [56]), 
            .I1(\edb_top_inst/la0/n1837 [11]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4528 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4529  (.I0(\edb_top_inst/edb_user_dr [57]), 
            .I1(\edb_top_inst/la0/n1837 [12]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4529 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4530  (.I0(\edb_top_inst/edb_user_dr [58]), 
            .I1(\edb_top_inst/la0/n1837 [13]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4530 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4531  (.I0(\edb_top_inst/edb_user_dr [59]), 
            .I1(\edb_top_inst/la0/n1837 [14]), .I2(\edb_top_inst/n2122 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4531 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4532  (.I0(\edb_top_inst/la0/n1837 [15]), 
            .I1(\edb_top_inst/la0/address_counter [15]), .I2(\edb_top_inst/n2134 ), 
            .O(\edb_top_inst/n2183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4532 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4533  (.I0(\edb_top_inst/n2183 ), .I1(\edb_top_inst/edb_user_dr [60]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4533 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4534  (.I0(\edb_top_inst/la0/n1837 [16]), 
            .I1(\edb_top_inst/la0/n1818 [1]), .I2(\edb_top_inst/n2134 ), 
            .O(\edb_top_inst/n2184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4534 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4535  (.I0(\edb_top_inst/n2184 ), .I1(\edb_top_inst/edb_user_dr [61]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4535 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4536  (.I0(\edb_top_inst/la0/n1818 [2]), .I1(\edb_top_inst/la0/n1837 [17]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4536 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4537  (.I0(\edb_top_inst/n2185 ), .I1(\edb_top_inst/edb_user_dr [62]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4537 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4538  (.I0(\edb_top_inst/la0/n1818 [3]), .I1(\edb_top_inst/la0/n1837 [18]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4538 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4539  (.I0(\edb_top_inst/n2186 ), .I1(\edb_top_inst/edb_user_dr [63]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4539 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4540  (.I0(\edb_top_inst/la0/n1818 [4]), .I1(\edb_top_inst/la0/n1837 [19]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4540 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4541  (.I0(\edb_top_inst/n2187 ), .I1(\edb_top_inst/edb_user_dr [64]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4541 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4542  (.I0(\edb_top_inst/la0/n1818 [5]), .I1(\edb_top_inst/la0/n1837 [20]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4542 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4543  (.I0(\edb_top_inst/n2188 ), .I1(\edb_top_inst/edb_user_dr [65]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4543 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4544  (.I0(\edb_top_inst/la0/n1818 [6]), .I1(\edb_top_inst/la0/n1837 [21]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4544 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4545  (.I0(\edb_top_inst/n2189 ), .I1(\edb_top_inst/edb_user_dr [66]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4545 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4546  (.I0(\edb_top_inst/la0/n1818 [7]), .I1(\edb_top_inst/la0/n1837 [22]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4546 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4547  (.I0(\edb_top_inst/n2190 ), .I1(\edb_top_inst/edb_user_dr [67]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4547 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4548  (.I0(\edb_top_inst/la0/n1818 [8]), .I1(\edb_top_inst/la0/n1837 [23]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4548 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4549  (.I0(\edb_top_inst/n2191 ), .I1(\edb_top_inst/edb_user_dr [68]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4549 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4550  (.I0(\edb_top_inst/la0/n1818 [9]), .I1(\edb_top_inst/la0/n1837 [24]), 
            .I2(\edb_top_inst/n2134 ), .O(\edb_top_inst/n2192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4550 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4551  (.I0(\edb_top_inst/n2192 ), .I1(\edb_top_inst/edb_user_dr [69]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_addr_counter [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4551 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4566  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/la0/n1984 [1]), 
            .O(\edb_top_inst/la0/n1998 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4566 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4567  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/la0/n1984 [2]), 
            .O(\edb_top_inst/la0/n1998 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4567 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4568  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/la0/n1984 [3]), 
            .O(\edb_top_inst/la0/n1998 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4568 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4569  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/la0/n1984 [4]), 
            .O(\edb_top_inst/la0/n1998 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4569 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4570  (.I0(\edb_top_inst/n2147 ), .I1(\edb_top_inst/la0/n1984 [5]), 
            .O(\edb_top_inst/la0/n1998 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4570 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4571  (.I0(\edb_top_inst/edb_user_dr [30]), 
            .I1(\edb_top_inst/la0/word_count [1]), .I2(\edb_top_inst/la0/word_count [0]), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4571 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__4572  (.I0(\edb_top_inst/la0/word_count [0]), 
            .I1(\edb_top_inst/la0/word_count [1]), .O(\edb_top_inst/n2200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4572 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4573  (.I0(\edb_top_inst/edb_user_dr [31]), 
            .I1(\edb_top_inst/la0/word_count [2]), .I2(\edb_top_inst/n2200 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4573 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4574  (.I0(\edb_top_inst/la0/word_count [2]), 
            .I1(\edb_top_inst/n2200 ), .I2(\edb_top_inst/la0/word_count [3]), 
            .O(\edb_top_inst/n2201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4574 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4575  (.I0(\edb_top_inst/n2201 ), .I1(\edb_top_inst/edb_user_dr [32]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4575 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4576  (.I0(\edb_top_inst/edb_user_dr [33]), 
            .I1(\edb_top_inst/la0/word_count [4]), .I2(\edb_top_inst/n2083 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4576 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4577  (.I0(\edb_top_inst/la0/word_count [4]), 
            .I1(\edb_top_inst/n2083 ), .O(\edb_top_inst/n2202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4577 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4578  (.I0(\edb_top_inst/edb_user_dr [34]), 
            .I1(\edb_top_inst/la0/word_count [5]), .I2(\edb_top_inst/n2202 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4578 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4579  (.I0(\edb_top_inst/la0/word_count [5]), 
            .I1(\edb_top_inst/n2202 ), .O(\edb_top_inst/n2203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4579 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4580  (.I0(\edb_top_inst/edb_user_dr [35]), 
            .I1(\edb_top_inst/la0/word_count [6]), .I2(\edb_top_inst/n2203 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4580 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4581  (.I0(\edb_top_inst/la0/word_count [6]), 
            .I1(\edb_top_inst/n2203 ), .O(\edb_top_inst/n2204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4581 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4582  (.I0(\edb_top_inst/edb_user_dr [36]), 
            .I1(\edb_top_inst/la0/word_count [7]), .I2(\edb_top_inst/n2204 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4582 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4583  (.I0(\edb_top_inst/n2083 ), .I1(\edb_top_inst/n2084 ), 
            .O(\edb_top_inst/n2205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4583 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4584  (.I0(\edb_top_inst/edb_user_dr [37]), 
            .I1(\edb_top_inst/la0/word_count [8]), .I2(\edb_top_inst/n2205 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4584 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4585  (.I0(\edb_top_inst/la0/word_count [8]), 
            .I1(\edb_top_inst/n2205 ), .O(\edb_top_inst/n2206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4585 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4586  (.I0(\edb_top_inst/edb_user_dr [38]), 
            .I1(\edb_top_inst/la0/word_count [9]), .I2(\edb_top_inst/n2206 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4586 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4587  (.I0(\edb_top_inst/la0/word_count [9]), 
            .I1(\edb_top_inst/n2206 ), .I2(\edb_top_inst/la0/word_count [10]), 
            .O(\edb_top_inst/n2207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4587 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4588  (.I0(\edb_top_inst/n2207 ), .I1(\edb_top_inst/edb_user_dr [39]), 
            .I2(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4588 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4589  (.I0(\edb_top_inst/n2205 ), .I1(\edb_top_inst/n2136 ), 
            .O(\edb_top_inst/n2208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4589 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4590  (.I0(\edb_top_inst/edb_user_dr [40]), 
            .I1(\edb_top_inst/la0/word_count [11]), .I2(\edb_top_inst/n2208 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4590 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4591  (.I0(\edb_top_inst/la0/word_count [11]), 
            .I1(\edb_top_inst/n2208 ), .O(\edb_top_inst/n2209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4591 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4592  (.I0(\edb_top_inst/edb_user_dr [41]), 
            .I1(\edb_top_inst/la0/word_count [12]), .I2(\edb_top_inst/n2209 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4592 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4593  (.I0(\edb_top_inst/la0/word_count [12]), 
            .I1(\edb_top_inst/n2209 ), .O(\edb_top_inst/n2210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4593 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4594  (.I0(\edb_top_inst/edb_user_dr [42]), 
            .I1(\edb_top_inst/la0/word_count [13]), .I2(\edb_top_inst/n2210 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4594 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4595  (.I0(\edb_top_inst/la0/word_count [12]), 
            .I1(\edb_top_inst/la0/word_count [13]), .I2(\edb_top_inst/n2209 ), 
            .O(\edb_top_inst/n2211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4595 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4596  (.I0(\edb_top_inst/edb_user_dr [43]), 
            .I1(\edb_top_inst/la0/word_count [14]), .I2(\edb_top_inst/n2211 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4596 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4597  (.I0(\edb_top_inst/la0/word_count [14]), 
            .I1(\edb_top_inst/n2211 ), .O(\edb_top_inst/n2212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4597 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4598  (.I0(\edb_top_inst/edb_user_dr [44]), 
            .I1(\edb_top_inst/la0/word_count [15]), .I2(\edb_top_inst/n2212 ), 
            .I3(\edb_top_inst/n2122 ), .O(\edb_top_inst/la0/data_to_word_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4598 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4599  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n2213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4599 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__4600  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4600 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4601  (.I0(\edb_top_inst/n2213 ), .I1(\edb_top_inst/la0/la_trig_mask [1]), 
            .I2(\edb_top_inst/n2214 ), .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4601 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__4602  (.I0(\edb_top_inst/la0/internal_register_select [1]), 
            .I1(\edb_top_inst/n2152 ), .I2(\edb_top_inst/n2153 ), .I3(\edb_top_inst/n2154 ), 
            .O(\edb_top_inst/n2216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4602 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4603  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/n2216 ), .O(\edb_top_inst/n2217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4603 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4604  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4604 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4605  (.I0(\edb_top_inst/n2218 ), .I1(\edb_top_inst/la0/skip_count [1]), 
            .I2(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4605 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4606  (.I0(\edb_top_inst/n2219 ), .I1(\edb_top_inst/n2215 ), 
            .I2(\edb_top_inst/la0/data_from_biu [1]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4606 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4607  (.I0(\edb_top_inst/n2220 ), .I1(\edb_top_inst/la0/data_out_shift_reg [2]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4607 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4608  (.I0(\edb_top_inst/la0/skip_count [2]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4608 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4609  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/n2222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4609 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4610  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .I2(\edb_top_inst/n2222 ), 
            .O(\edb_top_inst/n2223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4610 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4611  (.I0(\edb_top_inst/n2217 ), .I1(\edb_top_inst/n2221 ), 
            .I2(\edb_top_inst/n2223 ), .I3(\edb_top_inst/n2161 ), .O(\edb_top_inst/n2224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4611 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4612  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4612 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4613  (.I0(\edb_top_inst/la0/la_trig_mask [2]), 
            .I1(\edb_top_inst/n2225 ), .O(\edb_top_inst/n2226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4613 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4614  (.I0(\edb_top_inst/n2226 ), .I1(\edb_top_inst/n2224 ), 
            .I2(\edb_top_inst/la0/data_from_biu [2]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4614 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4615  (.I0(\edb_top_inst/n2227 ), .I1(\edb_top_inst/la0/data_out_shift_reg [3]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4615 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4616  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/la0/internal_register_select [0]), .I2(\edb_top_inst/n2216 ), 
            .O(\edb_top_inst/n2228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4616 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4617  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [3]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4617 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4618  (.I0(\edb_top_inst/la0/la_sample_cnt [0]), 
            .I1(\edb_top_inst/la0/la_trig_mask [3]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4618 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4619  (.I0(\edb_top_inst/n2230 ), .I1(\edb_top_inst/n2229 ), 
            .I2(\edb_top_inst/la0/data_from_biu [3]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4619 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4620  (.I0(\edb_top_inst/n2231 ), .I1(\edb_top_inst/la0/data_out_shift_reg [4]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4620 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4621  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/la0/internal_register_select [0]), .I2(\edb_top_inst/n2216 ), 
            .O(\edb_top_inst/n2232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4621 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__4622  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [4]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4622 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4623  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [4]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4623 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4624  (.I0(\edb_top_inst/n2234 ), .I1(\edb_top_inst/n2233 ), 
            .I2(\edb_top_inst/la0/data_from_biu [4]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4624 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4625  (.I0(\edb_top_inst/n2235 ), .I1(\edb_top_inst/la0/data_out_shift_reg [5]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4625 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4627  (.I0(\edb_top_inst/la0/la_sample_cnt [2]), 
            .I1(\edb_top_inst/la0/la_trig_mask [5]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4627 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4338  (.I0(\edb_top_inst/la0/crc_data_out [29]), 
            .I1(\edb_top_inst/edb_user_dr [79]), .I2(\edb_top_inst/la0/crc_data_out [30]), 
            .I3(\edb_top_inst/edb_user_dr [80]), .O(\edb_top_inst/n2055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4338 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4628  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [5]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2237 ), .O(\edb_top_inst/n2238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4628 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4629  (.I0(\edb_top_inst/n2238 ), .I1(\edb_top_inst/la0/data_from_biu [5]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4629 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4630  (.I0(\edb_top_inst/n2239 ), .I1(\edb_top_inst/la0/data_out_shift_reg [6]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4630 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4631  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/la0/la_sample_cnt [3]), 
            .I2(\edb_top_inst/la0/skip_count [6]), .I3(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4631 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4632  (.I0(\edb_top_inst/n2240 ), .I1(\edb_top_inst/la0/la_trig_mask [6]), 
            .I2(\edb_top_inst/n2225 ), .O(\edb_top_inst/n2241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4632 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4633  (.I0(\edb_top_inst/n2241 ), .I1(\edb_top_inst/la0/data_from_biu [6]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4633 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4634  (.I0(\edb_top_inst/n2242 ), .I1(\edb_top_inst/la0/data_out_shift_reg [7]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4634 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4635  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [7]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4635 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4636  (.I0(\edb_top_inst/la0/la_sample_cnt [4]), 
            .I1(\edb_top_inst/la0/la_trig_mask [7]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4636 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4637  (.I0(\edb_top_inst/n2244 ), .I1(\edb_top_inst/n2243 ), 
            .I2(\edb_top_inst/la0/data_from_biu [7]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4637 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4638  (.I0(\edb_top_inst/n2245 ), .I1(\edb_top_inst/la0/data_out_shift_reg [8]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4638 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4639  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [8]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4639 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4640  (.I0(\edb_top_inst/la0/la_sample_cnt [5]), 
            .I1(\edb_top_inst/la0/la_trig_mask [8]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4640 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4641  (.I0(\edb_top_inst/n2247 ), .I1(\edb_top_inst/n2246 ), 
            .I2(\edb_top_inst/la0/data_from_biu [8]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4641 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4642  (.I0(\edb_top_inst/n2248 ), .I1(\edb_top_inst/la0/data_out_shift_reg [9]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4642 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4643  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [9]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4643 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4644  (.I0(\edb_top_inst/la0/la_sample_cnt [6]), 
            .I1(\edb_top_inst/la0/la_trig_mask [9]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4644 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4645  (.I0(\edb_top_inst/n2250 ), .I1(\edb_top_inst/n2249 ), 
            .I2(\edb_top_inst/la0/data_from_biu [9]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4645 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4646  (.I0(\edb_top_inst/n2251 ), .I1(\edb_top_inst/la0/data_out_shift_reg [10]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4646 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4647  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [10]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4647 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4648  (.I0(\edb_top_inst/la0/la_sample_cnt [7]), 
            .I1(\edb_top_inst/la0/la_trig_mask [10]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4648 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4649  (.I0(\edb_top_inst/n2253 ), .I1(\edb_top_inst/n2252 ), 
            .I2(\edb_top_inst/la0/data_from_biu [10]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4649 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4650  (.I0(\edb_top_inst/n2254 ), .I1(\edb_top_inst/la0/data_out_shift_reg [11]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4650 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4651  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [11]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4651 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4652  (.I0(\edb_top_inst/la0/la_sample_cnt [8]), 
            .I1(\edb_top_inst/la0/la_trig_mask [11]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4652 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4653  (.I0(\edb_top_inst/n2256 ), .I1(\edb_top_inst/n2255 ), 
            .I2(\edb_top_inst/la0/data_from_biu [11]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4653 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4654  (.I0(\edb_top_inst/n2257 ), .I1(\edb_top_inst/la0/data_out_shift_reg [12]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4654 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4655  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [12]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4655 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4656  (.I0(\edb_top_inst/la0/la_sample_cnt [9]), 
            .I1(\edb_top_inst/la0/la_trig_mask [12]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4656 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4657  (.I0(\edb_top_inst/n2259 ), .I1(\edb_top_inst/n2258 ), 
            .I2(\edb_top_inst/la0/data_from_biu [12]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4657 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4658  (.I0(\edb_top_inst/n2260 ), .I1(\edb_top_inst/la0/data_out_shift_reg [13]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4658 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4659  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [13]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4659 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4660  (.I0(\edb_top_inst/la0/la_sample_cnt [10]), 
            .I1(\edb_top_inst/la0/la_trig_mask [13]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4660 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4661  (.I0(\edb_top_inst/n2262 ), .I1(\edb_top_inst/n2261 ), 
            .I2(\edb_top_inst/la0/data_from_biu [13]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4661 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4662  (.I0(\edb_top_inst/n2263 ), .I1(\edb_top_inst/la0/data_out_shift_reg [14]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4662 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4663  (.I0(\edb_top_inst/la0/skip_count [14]), 
            .I1(\edb_top_inst/n2156 ), .I2(\edb_top_inst/n2218 ), .O(\edb_top_inst/n2264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4663 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4664  (.I0(\edb_top_inst/la0/la_trig_mask [14]), 
            .I1(\edb_top_inst/la0/data_from_biu [14]), .I2(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4664 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4665  (.I0(\edb_top_inst/n2264 ), .I1(\edb_top_inst/n2265 ), 
            .I2(\edb_top_inst/n2225 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5cc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4665 .LUTMASK = 16'hc5cc;
    EFX_LUT4 \edb_top_inst/LUT__4666  (.I0(\edb_top_inst/n2266 ), .I1(\edb_top_inst/la0/data_out_shift_reg [15]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4666 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4667  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4667 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4668  (.I0(\edb_top_inst/la0/skip_count [15]), 
            .I1(\edb_top_inst/n2156 ), .I2(\edb_top_inst/n2267 ), .O(\edb_top_inst/n2268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4668 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4669  (.I0(\edb_top_inst/la0/la_trig_mask [15]), 
            .I1(\edb_top_inst/la0/data_from_biu [15]), .I2(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4669 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4670  (.I0(\edb_top_inst/n2268 ), .I1(\edb_top_inst/n2269 ), 
            .I2(\edb_top_inst/n2225 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5cc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4670 .LUTMASK = 16'hc5cc;
    EFX_LUT4 \edb_top_inst/LUT__4671  (.I0(\edb_top_inst/n2270 ), .I1(\edb_top_inst/la0/data_out_shift_reg [16]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4671 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4672  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [16]), 
            .I2(\edb_top_inst/la0/la_trig_mask [16]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4672 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4673  (.I0(\edb_top_inst/n2271 ), .I1(\edb_top_inst/la0/data_from_biu [16]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4673 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4674  (.I0(\edb_top_inst/n2272 ), .I1(\edb_top_inst/la0/data_out_shift_reg [17]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4674 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4675  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4675 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4676  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [17]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2273 ), .O(\edb_top_inst/n2274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4676 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4677  (.I0(\edb_top_inst/n2274 ), .I1(\edb_top_inst/la0/data_from_biu [17]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4677 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4678  (.I0(\edb_top_inst/n2275 ), .I1(\edb_top_inst/la0/data_out_shift_reg [18]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4678 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4679  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [18]), 
            .I2(\edb_top_inst/la0/la_trig_mask [18]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4679 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4680  (.I0(\edb_top_inst/n2276 ), .I1(\edb_top_inst/la0/data_from_biu [18]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4680 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4681  (.I0(\edb_top_inst/n2277 ), .I1(\edb_top_inst/la0/data_out_shift_reg [19]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4681 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4682  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [19]), 
            .I2(\edb_top_inst/la0/la_trig_mask [19]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4682 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4683  (.I0(\edb_top_inst/n2278 ), .I1(\edb_top_inst/la0/data_from_biu [19]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4683 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4684  (.I0(\edb_top_inst/n2279 ), .I1(\edb_top_inst/la0/data_out_shift_reg [20]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4684 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4685  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [20]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4685 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4686  (.I0(\edb_top_inst/la0/la_trig_mask [20]), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4686 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4687  (.I0(\edb_top_inst/n2281 ), .I1(\edb_top_inst/n2280 ), 
            .I2(\edb_top_inst/la0/data_from_biu [20]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4687 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4688  (.I0(\edb_top_inst/n2282 ), .I1(\edb_top_inst/la0/data_out_shift_reg [21]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4688 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4689  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [21]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4689 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4690  (.I0(\edb_top_inst/la0/la_trig_mask [21]), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4690 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4691  (.I0(\edb_top_inst/n2284 ), .I1(\edb_top_inst/n2283 ), 
            .I2(\edb_top_inst/la0/data_from_biu [21]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4691 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4692  (.I0(\edb_top_inst/n2285 ), .I1(\edb_top_inst/la0/data_out_shift_reg [22]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4692 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4693  (.I0(\edb_top_inst/la0/la_trig_mask [22]), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4693 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4694  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [22]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2286 ), .O(\edb_top_inst/n2287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4694 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4695  (.I0(\edb_top_inst/n2287 ), .I1(\edb_top_inst/la0/data_from_biu [22]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4695 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4696  (.I0(\edb_top_inst/n2288 ), .I1(\edb_top_inst/la0/data_out_shift_reg [23]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4696 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4697  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_trig_mask [23]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4697 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4698  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [23]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2289 ), .O(\edb_top_inst/n2290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4698 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4699  (.I0(\edb_top_inst/n2290 ), .I1(\edb_top_inst/la0/data_from_biu [23]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4699 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4700  (.I0(\edb_top_inst/n2291 ), .I1(\edb_top_inst/la0/data_out_shift_reg [24]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4700 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4701  (.I0(\edb_top_inst/la0/la_trig_pos [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [24]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4701 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4702  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [24]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2292 ), .O(\edb_top_inst/n2293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4702 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4703  (.I0(\edb_top_inst/n2293 ), .I1(\edb_top_inst/la0/data_from_biu [24]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4703 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4704  (.I0(\edb_top_inst/n2294 ), .I1(\edb_top_inst/la0/data_out_shift_reg [25]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4704 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4705  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [25]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4705 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4706  (.I0(\edb_top_inst/la0/la_trig_pos [2]), 
            .I1(\edb_top_inst/la0/la_trig_mask [25]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4706 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4707  (.I0(\edb_top_inst/n2296 ), .I1(\edb_top_inst/n2295 ), 
            .I2(\edb_top_inst/la0/data_from_biu [25]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4707 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4708  (.I0(\edb_top_inst/n2297 ), .I1(\edb_top_inst/la0/data_out_shift_reg [26]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4708 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4709  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [26]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4709 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4710  (.I0(\edb_top_inst/la0/la_trig_pos [3]), 
            .I1(\edb_top_inst/la0/la_trig_mask [26]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4710 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4711  (.I0(\edb_top_inst/n2299 ), .I1(\edb_top_inst/n2298 ), 
            .I2(\edb_top_inst/la0/data_from_biu [26]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4711 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4712  (.I0(\edb_top_inst/n2300 ), .I1(\edb_top_inst/la0/data_out_shift_reg [27]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4712 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4713  (.I0(\edb_top_inst/la0/la_trig_pos [4]), 
            .I1(\edb_top_inst/la0/la_trig_mask [27]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4713 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4714  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [27]), 
            .I2(\edb_top_inst/n2159 ), .I3(\edb_top_inst/n2218 ), .O(\edb_top_inst/n2302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4714 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__4715  (.I0(\edb_top_inst/n2302 ), .I1(\edb_top_inst/n2301 ), 
            .I2(\edb_top_inst/la0/data_from_biu [27]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4715 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4716  (.I0(\edb_top_inst/n2303 ), .I1(\edb_top_inst/la0/data_out_shift_reg [28]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4716 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4717  (.I0(\edb_top_inst/la0/la_trig_pos [5]), 
            .I1(\edb_top_inst/la0/la_trig_mask [28]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4717 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4718  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [28]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2304 ), .O(\edb_top_inst/n2305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4718 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4719  (.I0(\edb_top_inst/n2305 ), .I1(\edb_top_inst/la0/data_from_biu [28]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4719 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4720  (.I0(\edb_top_inst/n2306 ), .I1(\edb_top_inst/la0/data_out_shift_reg [29]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4720 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4721  (.I0(\edb_top_inst/la0/la_trig_pos [6]), 
            .I1(\edb_top_inst/la0/la_trig_mask [29]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4721 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4722  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [29]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2307 ), .O(\edb_top_inst/n2308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4722 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4723  (.I0(\edb_top_inst/n2308 ), .I1(\edb_top_inst/la0/data_from_biu [29]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4723 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4724  (.I0(\edb_top_inst/n2309 ), .I1(\edb_top_inst/la0/data_out_shift_reg [30]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4724 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4725  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [30]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4725 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4726  (.I0(\edb_top_inst/la0/la_trig_pos [7]), 
            .I1(\edb_top_inst/la0/la_trig_mask [30]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4726 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4727  (.I0(\edb_top_inst/n2311 ), .I1(\edb_top_inst/n2310 ), 
            .I2(\edb_top_inst/la0/data_from_biu [30]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4727 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4728  (.I0(\edb_top_inst/n2312 ), .I1(\edb_top_inst/la0/data_out_shift_reg [31]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4728 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4729  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [31]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4729 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4730  (.I0(\edb_top_inst/la0/la_trig_pos [8]), 
            .I1(\edb_top_inst/la0/la_trig_mask [31]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4730 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4731  (.I0(\edb_top_inst/n2314 ), .I1(\edb_top_inst/n2313 ), 
            .I2(\edb_top_inst/la0/data_from_biu [31]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4731 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4732  (.I0(\edb_top_inst/n2315 ), .I1(\edb_top_inst/la0/data_out_shift_reg [32]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4732 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4733  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/la0/la_trig_pos [9]), 
            .I2(\edb_top_inst/la0/skip_count [32]), .I3(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4733 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4734  (.I0(\edb_top_inst/n2316 ), .I1(\edb_top_inst/la0/la_trig_mask [32]), 
            .I2(\edb_top_inst/n2225 ), .O(\edb_top_inst/n2317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4734 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4735  (.I0(\edb_top_inst/n2317 ), .I1(\edb_top_inst/la0/data_from_biu [32]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4735 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4736  (.I0(\edb_top_inst/n2318 ), .I1(\edb_top_inst/la0/data_out_shift_reg [33]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4736 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4737  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/la0/la_trig_pos [10]), 
            .I2(\edb_top_inst/la0/skip_count [33]), .I3(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4737 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4738  (.I0(\edb_top_inst/n2319 ), .I1(\edb_top_inst/la0/la_trig_mask [33]), 
            .I2(\edb_top_inst/n2225 ), .O(\edb_top_inst/n2320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4738 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4739  (.I0(\edb_top_inst/n2320 ), .I1(\edb_top_inst/la0/data_from_biu [33]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4739 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4740  (.I0(\edb_top_inst/n2321 ), .I1(\edb_top_inst/la0/data_out_shift_reg [34]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4740 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4741  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [34]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4741 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4742  (.I0(\edb_top_inst/la0/la_trig_pos [11]), 
            .I1(\edb_top_inst/la0/la_trig_mask [34]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4742 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4743  (.I0(\edb_top_inst/n2323 ), .I1(\edb_top_inst/n2322 ), 
            .I2(\edb_top_inst/la0/data_from_biu [34]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4743 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4744  (.I0(\edb_top_inst/n2324 ), .I1(\edb_top_inst/la0/data_out_shift_reg [35]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4744 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4745  (.I0(\edb_top_inst/la0/la_trig_pos [12]), 
            .I1(\edb_top_inst/la0/la_trig_mask [35]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4745 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4746  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [35]), 
            .I2(\edb_top_inst/n2217 ), .I3(\edb_top_inst/n2325 ), .O(\edb_top_inst/n2326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4746 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4747  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/la0/data_from_biu [35]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4747 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4748  (.I0(\edb_top_inst/n2327 ), .I1(\edb_top_inst/la0/data_out_shift_reg [36]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4748 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4749  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [36]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4749 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4750  (.I0(\edb_top_inst/la0/la_trig_pos [13]), 
            .I1(\edb_top_inst/la0/la_trig_mask [36]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4750 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4751  (.I0(\edb_top_inst/n2329 ), .I1(\edb_top_inst/n2328 ), 
            .I2(\edb_top_inst/la0/data_from_biu [36]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4751 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4752  (.I0(\edb_top_inst/n2330 ), .I1(\edb_top_inst/la0/data_out_shift_reg [37]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4752 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4753  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [37]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4753 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4754  (.I0(\edb_top_inst/la0/la_trig_pos [14]), 
            .I1(\edb_top_inst/la0/la_trig_mask [37]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4754 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4755  (.I0(\edb_top_inst/n2332 ), .I1(\edb_top_inst/n2331 ), 
            .I2(\edb_top_inst/la0/data_from_biu [37]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4755 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4756  (.I0(\edb_top_inst/n2333 ), .I1(\edb_top_inst/la0/data_out_shift_reg [38]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4756 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4757  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [38]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4757 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4758  (.I0(\edb_top_inst/la0/la_trig_pos [15]), 
            .I1(\edb_top_inst/la0/la_trig_mask [38]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4758 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4759  (.I0(\edb_top_inst/n2335 ), .I1(\edb_top_inst/n2334 ), 
            .I2(\edb_top_inst/la0/data_from_biu [38]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4759 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4760  (.I0(\edb_top_inst/n2336 ), .I1(\edb_top_inst/la0/data_out_shift_reg [39]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4760 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4761  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/la0/la_trig_pos [16]), 
            .I2(\edb_top_inst/la0/skip_count [39]), .I3(\edb_top_inst/n2156 ), 
            .O(\edb_top_inst/n2337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4761 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4762  (.I0(\edb_top_inst/n2337 ), .I1(\edb_top_inst/la0/la_trig_mask [39]), 
            .I2(\edb_top_inst/n2225 ), .O(\edb_top_inst/n2338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4762 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4763  (.I0(\edb_top_inst/n2338 ), .I1(\edb_top_inst/la0/data_from_biu [39]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4763 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4764  (.I0(\edb_top_inst/n2339 ), .I1(\edb_top_inst/la0/data_out_shift_reg [40]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4764 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4765  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [40]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4765 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4766  (.I0(\edb_top_inst/la0/la_trig_mask [40]), 
            .I1(\edb_top_inst/la0/la_trig_pattern [0]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4766 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4767  (.I0(\edb_top_inst/n2341 ), .I1(\edb_top_inst/n2340 ), 
            .I2(\edb_top_inst/la0/data_from_biu [40]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4767 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4768  (.I0(\edb_top_inst/n2342 ), .I1(\edb_top_inst/la0/data_out_shift_reg [41]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4768 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4769  (.I0(\edb_top_inst/la0/la_trig_mask [41]), 
            .I1(\edb_top_inst/la0/la_trig_pattern [1]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4769 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4770  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [41]), 
            .I2(\edb_top_inst/n2159 ), .I3(\edb_top_inst/n2218 ), .O(\edb_top_inst/n2344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4770 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__4771  (.I0(\edb_top_inst/n2344 ), .I1(\edb_top_inst/n2343 ), 
            .I2(\edb_top_inst/la0/data_from_biu [41]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4771 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4772  (.I0(\edb_top_inst/n2345 ), .I1(\edb_top_inst/la0/data_out_shift_reg [42]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4772 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4773  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [42]), 
            .I2(\edb_top_inst/n2232 ), .O(\edb_top_inst/n2346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4773 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4774  (.I0(\edb_top_inst/la0/la_trig_mask [42]), 
            .I1(\edb_top_inst/la0/la_capture_pattern [0]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2347 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4774 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4775  (.I0(\edb_top_inst/n2347 ), .I1(\edb_top_inst/n2346 ), 
            .I2(\edb_top_inst/la0/data_from_biu [42]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4775 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4776  (.I0(\edb_top_inst/n2348 ), .I1(\edb_top_inst/la0/data_out_shift_reg [43]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4776 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4777  (.I0(\edb_top_inst/n2214 ), .I1(\edb_top_inst/la0/skip_count [43]), 
            .I2(\edb_top_inst/n2228 ), .O(\edb_top_inst/n2349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4777 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4778  (.I0(\edb_top_inst/la0/la_trig_mask [43]), 
            .I1(\edb_top_inst/la0/la_capture_pattern [1]), .I2(\edb_top_inst/n2214 ), 
            .I3(\edb_top_inst/n2159 ), .O(\edb_top_inst/n2350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4778 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__4779  (.I0(\edb_top_inst/n2350 ), .I1(\edb_top_inst/n2349 ), 
            .I2(\edb_top_inst/la0/data_from_biu [43]), .I3(\edb_top_inst/n2164 ), 
            .O(\edb_top_inst/n2351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4779 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4780  (.I0(\edb_top_inst/n2351 ), .I1(\edb_top_inst/la0/data_out_shift_reg [44]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4780 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4781  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [44]), 
            .I2(\edb_top_inst/la0/la_trig_mask [44]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4781 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4782  (.I0(\edb_top_inst/n2352 ), .I1(\edb_top_inst/la0/data_from_biu [44]), 
            .I2(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2353 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4782 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__4783  (.I0(\edb_top_inst/n2353 ), .I1(\edb_top_inst/la0/data_out_shift_reg [45]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4783 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4784  (.I0(\edb_top_inst/la0/skip_count [45]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4784 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4785  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [45]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2354 ), .O(\edb_top_inst/n2355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4785 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4786  (.I0(\edb_top_inst/n2355 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [46]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4786 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4787  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [46]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4787 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4788  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [46]), 
            .I2(\edb_top_inst/n2356 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4788 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4789  (.I0(\edb_top_inst/n2357 ), .I1(\edb_top_inst/la0/data_out_shift_reg [47]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4789 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4790  (.I0(\edb_top_inst/la0/skip_count [47]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4790 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4791  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [47]), 
            .I2(\edb_top_inst/n2218 ), .I3(\edb_top_inst/n2358 ), .O(\edb_top_inst/n2359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4791 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4792  (.I0(\edb_top_inst/n2359 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [48]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4792 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4793  (.I0(\edb_top_inst/la0/skip_count [48]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4793 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4794  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [48]), 
            .I2(\edb_top_inst/n2218 ), .I3(\edb_top_inst/n2360 ), .O(\edb_top_inst/n2361 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4794 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4795  (.I0(\edb_top_inst/n2361 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [49]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4795 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4796  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [49]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4796 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4797  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [49]), 
            .I2(\edb_top_inst/n2362 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4797 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4798  (.I0(\edb_top_inst/n2363 ), .I1(\edb_top_inst/la0/data_out_shift_reg [50]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4798 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4799  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [50]), 
            .I2(\edb_top_inst/la0/la_trig_mask [50]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4799 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4800  (.I0(\edb_top_inst/n2364 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [51]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4800 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4801  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [51]), 
            .I2(\edb_top_inst/la0/la_trig_mask [51]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2365 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4801 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4802  (.I0(\edb_top_inst/n2365 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [52]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4802 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4803  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4803 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4804  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [52]), 
            .I2(\edb_top_inst/n2218 ), .I3(\edb_top_inst/n2366 ), .O(\edb_top_inst/n2367 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4804 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4805  (.I0(\edb_top_inst/n2367 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [53]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4805 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4806  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [53]), 
            .I2(\edb_top_inst/la0/la_trig_mask [53]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4806 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4807  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [54]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4807 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4808  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [54]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4808 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4809  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [54]), 
            .I2(\edb_top_inst/n2369 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4809 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4810  (.I0(\edb_top_inst/n2370 ), .I1(\edb_top_inst/la0/data_out_shift_reg [55]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4810 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4811  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4811 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4812  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [55]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2371 ), .O(\edb_top_inst/n2372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4812 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4813  (.I0(\edb_top_inst/n2372 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [56]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4813 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4814  (.I0(\edb_top_inst/la0/skip_count [56]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4814 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4815  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [56]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2373 ), .O(\edb_top_inst/n2374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4815 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4816  (.I0(\edb_top_inst/n2374 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [57]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4816 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4817  (.I0(\edb_top_inst/la0/skip_count [57]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4817 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4818  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [57]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2375 ), .O(\edb_top_inst/n2376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4818 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4819  (.I0(\edb_top_inst/n2376 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [58]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4819 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4820  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4820 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4821  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [58]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2377 ), .O(\edb_top_inst/n2378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4821 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4822  (.I0(\edb_top_inst/n2378 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [59]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4822 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4823  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [59]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4823 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4824  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [59]), 
            .I2(\edb_top_inst/n2379 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4824 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4825  (.I0(\edb_top_inst/n2380 ), .I1(\edb_top_inst/la0/data_out_shift_reg [60]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4825 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4826  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [60]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4826 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4827  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [60]), 
            .I2(\edb_top_inst/n2381 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4827 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4828  (.I0(\edb_top_inst/n2382 ), .I1(\edb_top_inst/la0/data_out_shift_reg [61]), 
            .I2(\edb_top_inst/n2168 ), .O(\edb_top_inst/la0/n2217 [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4828 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4829  (.I0(\edb_top_inst/la0/skip_count [61]), 
            .I1(\edb_top_inst/n2156 ), .O(\edb_top_inst/n2383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4829 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4830  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [61]), 
            .I2(\edb_top_inst/n2267 ), .I3(\edb_top_inst/n2383 ), .O(\edb_top_inst/n2384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4830 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4831  (.I0(\edb_top_inst/n2384 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [62]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4831 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4832  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [62]), 
            .I2(\edb_top_inst/la0/la_trig_mask [62]), .I3(\edb_top_inst/n2225 ), 
            .O(\edb_top_inst/n2385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4832 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4833  (.I0(\edb_top_inst/n2385 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [63]), .I3(\edb_top_inst/n2168 ), 
            .O(\edb_top_inst/la0/n2217 [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4833 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__4834  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/la0/skip_count [63]), 
            .I2(\edb_top_inst/n2217 ), .O(\edb_top_inst/n2386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4834 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4835  (.I0(\edb_top_inst/n2225 ), .I1(\edb_top_inst/la0/la_trig_mask [63]), 
            .I2(\edb_top_inst/n2386 ), .I3(\edb_top_inst/n2164 ), .O(\edb_top_inst/n2387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4835 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4836  (.I0(\edb_top_inst/n2168 ), .I1(\edb_top_inst/n2387 ), 
            .O(\edb_top_inst/la0/n2217 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4836 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4837  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/n2101 ), .I2(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n2388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4837 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4838  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n2389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f57, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4838 .LUTMASK = 16'h0f57;
    EFX_LUT4 \edb_top_inst/LUT__4839  (.I0(\edb_top_inst/n2087 ), .I1(\edb_top_inst/n2079 ), 
            .I2(\edb_top_inst/n2389 ), .I3(\edb_top_inst/la0/module_state [1]), 
            .O(\edb_top_inst/n2390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4839 .LUTMASK = 16'h0bbb;
    EFX_LUT4 \edb_top_inst/LUT__4840  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/n2079 ), .I2(\edb_top_inst/n2108 ), .O(\edb_top_inst/n2391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4840 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4841  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/n2390 ), .I2(\edb_top_inst/n2388 ), .I3(\edb_top_inst/n2391 ), 
            .O(\edb_top_inst/la0/module_next_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4841 .LUTMASK = 16'hff01;
    EFX_LUT4 \edb_top_inst/LUT__4842  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/n2150 ), .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n2088 ), 
            .O(\edb_top_inst/n2392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4842 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4843  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/n2094 ), .I2(\edb_top_inst/n2150 ), .I3(\edb_top_inst/n2087 ), 
            .O(\edb_top_inst/n2393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4843 .LUTMASK = 16'he800;
    EFX_LUT4 \edb_top_inst/LUT__4844  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n2087 ), 
            .I2(\edb_top_inst/n2144 ), .O(\edb_top_inst/n2394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4844 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4845  (.I0(\edb_top_inst/n2393 ), .I1(\edb_top_inst/n2392 ), 
            .I2(\edb_top_inst/n2140 ), .I3(\edb_top_inst/n2394 ), .O(\edb_top_inst/la0/module_next_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4845 .LUTMASK = 16'hfff4;
    EFX_LUT4 \edb_top_inst/LUT__4846  (.I0(\edb_top_inst/la0/crc_data_out [1]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4846 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4847  (.I0(\edb_top_inst/n2079 ), .I1(\edb_top_inst/n2097 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n2149 ), 
            .O(\edb_top_inst/ceg_net11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4847 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4848  (.I0(\edb_top_inst/la0/crc_data_out [2]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4848 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4849  (.I0(\edb_top_inst/la0/crc_data_out [3]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4849 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4850  (.I0(\edb_top_inst/la0/crc_data_out [4]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4850 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4851  (.I0(\edb_top_inst/la0/crc_data_out [5]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4851 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4852  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg [0]), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/la0/crc_data_out [0]), 
            .O(\edb_top_inst/n2395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4852 .LUTMASK = 16'h53ac;
    EFX_LUT4 \edb_top_inst/LUT__4853  (.I0(\edb_top_inst/n2079 ), .I1(\edb_top_inst/n2395 ), 
            .I2(\edb_top_inst/n2088 ), .O(\edb_top_inst/n2396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4853 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4854  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/n2396 ), .O(\edb_top_inst/n2397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4854 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4855  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [6]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4855 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4856  (.I0(\edb_top_inst/la0/crc_data_out [7]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4856 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4857  (.I0(\edb_top_inst/la0/crc_data_out [8]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4857 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4858  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [9]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4858 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4859  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [10]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4859 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4860  (.I0(\edb_top_inst/la0/crc_data_out [11]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4860 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4861  (.I0(\edb_top_inst/la0/crc_data_out [12]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4861 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4862  (.I0(\edb_top_inst/la0/crc_data_out [13]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4862 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4863  (.I0(\edb_top_inst/la0/crc_data_out [14]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4863 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4864  (.I0(\edb_top_inst/la0/crc_data_out [15]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4864 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4865  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [16]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4865 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4866  (.I0(\edb_top_inst/la0/crc_data_out [17]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4866 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4867  (.I0(\edb_top_inst/la0/crc_data_out [18]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4867 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4868  (.I0(\edb_top_inst/la0/crc_data_out [19]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4868 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4869  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [20]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4869 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4870  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [21]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4870 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4871  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [22]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4871 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4872  (.I0(\edb_top_inst/la0/crc_data_out [23]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4872 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4873  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [24]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4873 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4874  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [25]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4874 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4875  (.I0(\edb_top_inst/la0/crc_data_out [26]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4875 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4876  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [27]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4876 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4877  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [28]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4877 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4878  (.I0(\edb_top_inst/la0/crc_data_out [29]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4878 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4879  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [30]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4879 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4880  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [31]), .I2(\edb_top_inst/n2397 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4880 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4881  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n2397 ), .O(\edb_top_inst/la0/axi_crc_i/n118 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4881 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4882  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4882 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4883  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4883 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4884  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4884 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4885  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4885 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4886  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4886 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4887  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2398 ), .O(\edb_top_inst/n2399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4887 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4888  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4888 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4889  (.I0(\edb_top_inst/n2400 ), .I1(\edb_top_inst/n2399 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4889 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4890  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4890 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4891  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4891 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4892  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), .O(\edb_top_inst/n2401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4892 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4893  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n2401 ), .O(\edb_top_inst/n2402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4893 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4894  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I2(\edb_top_inst/n2402 ), .O(\edb_top_inst/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4894 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4895  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I2(\edb_top_inst/n2403 ), .O(\edb_top_inst/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4895 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4896  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/n2404 ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4896 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__4897  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I2(\edb_top_inst/n2405 ), .O(\edb_top_inst/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4897 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4898  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I2(\edb_top_inst/n2406 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4898 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4899  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4899 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4900  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4900 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4901  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4901 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4902  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4902 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4903  (.I0(\edb_top_inst/n2407 ), .I1(\edb_top_inst/n2408 ), 
            .I2(\edb_top_inst/n2409 ), .I3(\edb_top_inst/n2410 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4903 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4904  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4904 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4905  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4905 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4906  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4906 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4907  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5]), 
            .O(\edb_top_inst/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4907 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4908  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4908 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4909  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7]), 
            .O(\edb_top_inst/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4909 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4910  (.I0(\edb_top_inst/n2413 ), .I1(\edb_top_inst/n2414 ), 
            .I2(\edb_top_inst/n2415 ), .I3(\edb_top_inst/n2416 ), .O(\edb_top_inst/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4910 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4911  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/n2412 ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/n2417 ), .O(\edb_top_inst/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2f75, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4911 .LUTMASK = 16'h2f75;
    EFX_LUT4 \edb_top_inst/LUT__4912  (.I0(\edb_top_inst/n2418 ), .I1(\edb_top_inst/n2411 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4912 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4913  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4913 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4914  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4914 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4915  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4915 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4916  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4916 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4917  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4917 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4918  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4918 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4919  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4919 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4920  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4920 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4921  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4921 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4922  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4922 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4923  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4923 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4924  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4924 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4925  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4925 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4926  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4926 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4927  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4927 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4928  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4928 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4929  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4929 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4930  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4930 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4931  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4931 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4932  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/n2419 ), .O(\edb_top_inst/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4932 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4933  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4933 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4934  (.I0(\edb_top_inst/n2421 ), .I1(\edb_top_inst/n2420 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4934 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4935  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4935 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4936  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4936 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4937  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4937 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4938  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4938 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4939  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4939 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4940  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2422 ), .O(\edb_top_inst/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4940 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4941  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4941 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4942  (.I0(\edb_top_inst/n2424 ), .I1(\edb_top_inst/n2423 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4942 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4943  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4943 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4944  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4944 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4945  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4945 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4946  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4946 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4947  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4947 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4948  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/n2425 ), .O(\edb_top_inst/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4948 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4949  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4949 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4950  (.I0(\edb_top_inst/n2427 ), .I1(\edb_top_inst/n2426 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4950 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4955  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4955 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4956  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2428 ), .O(\edb_top_inst/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4956 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4957  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4957 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4958  (.I0(\edb_top_inst/n2430 ), .I1(\edb_top_inst/n2429 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4958 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4959  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4959 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4960  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4960 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4961  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4961 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4962  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4962 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4963  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4963 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4964  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2431 ), .O(\edb_top_inst/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4964 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4965  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4965 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4966  (.I0(\edb_top_inst/n2433 ), .I1(\edb_top_inst/n2432 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4966 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4967  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4967 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4968  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4968 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4969  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), .O(\edb_top_inst/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4969 .LUTMASK = 16'hefef;
    EFX_LUT4 \edb_top_inst/LUT__4970  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/n2434 ), .O(\edb_top_inst/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4970 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4971  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/n2435 ), .O(\edb_top_inst/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4971 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4972  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I2(\edb_top_inst/n2436 ), .O(\edb_top_inst/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4972 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4973  (.I0(\edb_top_inst/n2437 ), .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdddd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4973 .LUTMASK = 16'hdddd;
    EFX_LUT4 \edb_top_inst/LUT__4974  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I1(\edb_top_inst/n2438 ), .O(\edb_top_inst/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4974 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4975  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I1(\edb_top_inst/n2439 ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4975 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4976  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4976 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4977  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4977 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4978  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4978 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4979  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4979 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4980  (.I0(\edb_top_inst/n2440 ), .I1(\edb_top_inst/n2441 ), 
            .I2(\edb_top_inst/n2442 ), .I3(\edb_top_inst/n2443 ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4980 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4981  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4981 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__4982  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4982 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4983  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5]), 
            .O(\edb_top_inst/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4983 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4984  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4984 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4985  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7]), 
            .O(\edb_top_inst/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4985 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4986  (.I0(\edb_top_inst/n2445 ), .I1(\edb_top_inst/n2446 ), 
            .I2(\edb_top_inst/n2447 ), .I3(\edb_top_inst/n2448 ), .O(\edb_top_inst/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4986 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4987  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I3(\edb_top_inst/n2449 ), .O(\edb_top_inst/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4987 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4988  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4988 .LUTMASK = 16'h1ff3;
    EFX_LUT4 \edb_top_inst/LUT__4989  (.I0(\edb_top_inst/n2444 ), .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/n2450 ), .I3(\edb_top_inst/n2451 ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4989 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4990  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4990 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4991  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4991 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4992  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4992 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4993  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4993 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4994  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4994 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4995  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4995 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4996  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n32 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4996 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4997  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4997 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4998  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4998 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4999  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4999 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5000  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5000 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5001  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5001 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5002  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5002 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5003  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n14 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5003 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5004  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5004 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5005  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5005 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5006  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), .O(\edb_top_inst/n2452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5006 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__5007  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n2452 ), .O(\edb_top_inst/n2453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5007 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__5008  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I2(\edb_top_inst/n2453 ), .O(\edb_top_inst/n2454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5008 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__5009  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I2(\edb_top_inst/n2454 ), .O(\edb_top_inst/n2455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5009 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__5010  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/n2455 ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/n2456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5010 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__5011  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I2(\edb_top_inst/n2456 ), .O(\edb_top_inst/n2457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5011 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__5012  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I2(\edb_top_inst/n2457 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5012 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__5013  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/n2458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5013 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5014  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/n2459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5014 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5015  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5015 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5016  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/n2461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5016 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5017  (.I0(\edb_top_inst/n2458 ), .I1(\edb_top_inst/n2459 ), 
            .I2(\edb_top_inst/n2460 ), .I3(\edb_top_inst/n2461 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5017 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__5018  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/n2462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5018 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__5019  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5019 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5020  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5]), 
            .O(\edb_top_inst/n2464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5020 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5021  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5021 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5022  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7]), 
            .O(\edb_top_inst/n2466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5022 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5023  (.I0(\edb_top_inst/n2463 ), .I1(\edb_top_inst/n2464 ), 
            .I2(\edb_top_inst/n2465 ), .I3(\edb_top_inst/n2466 ), .O(\edb_top_inst/n2467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5023 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5024  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I3(\edb_top_inst/n2467 ), .O(\edb_top_inst/n2468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5024 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__5025  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5025 .LUTMASK = 16'h1ff3;
    EFX_LUT4 \edb_top_inst/LUT__5026  (.I0(\edb_top_inst/n2462 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/n2468 ), .I3(\edb_top_inst/n2469 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5026 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__5027  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5027 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5028  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5028 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5029  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5029 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5030  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5030 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5031  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5031 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5032  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5032 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5033  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n32 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5033 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5034  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5034 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5035  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5035 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5036  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5036 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5037  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5037 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5038  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5038 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5039  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5039 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5040  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n14 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5040 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5041  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5041 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5042  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5042 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5043  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [0]), .O(\edb_top_inst/n2470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5043 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__5044  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [3]), .O(\edb_top_inst/n2471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5044 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__5045  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [3]), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5045 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5046  (.I0(\edb_top_inst/n2471 ), .I1(\edb_top_inst/n2470 ), 
            .I2(\edb_top_inst/n2472 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5046 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__5047  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [1]), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5047 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5048  (.I0(\edb_top_inst/n2472 ), .I1(\edb_top_inst/n2473 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5048 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__5049  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5049 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__5050  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/n2474 ), .O(\edb_top_inst/n2475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8c3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5050 .LUTMASK = 16'ha8c3;
    EFX_LUT4 \edb_top_inst/LUT__5051  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5051 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5052  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5052 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5053  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/n2476 ), .I3(\edb_top_inst/n2477 ), .O(\edb_top_inst/n2478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5053 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__5054  (.I0(\edb_top_inst/n2478 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n2475 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5054 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__5055  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5055 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5056  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5056 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5057  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5057 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5058  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5058 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5059  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5059 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5060  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n10 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5060 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5061  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5061 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5062  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5062 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5063  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [0]), .O(\edb_top_inst/n2479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5063 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__5064  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [3]), .O(\edb_top_inst/n2480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5064 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__5065  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [3]), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5065 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5066  (.I0(\edb_top_inst/n2480 ), .I1(\edb_top_inst/n2479 ), 
            .I2(\edb_top_inst/n2481 ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5066 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__5067  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [1]), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5067 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5068  (.I0(\edb_top_inst/n2481 ), .I1(\edb_top_inst/n2482 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/equal_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5068 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__5069  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5069 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__5070  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n2483 ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he83f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5070 .LUTMASK = 16'he83f;
    EFX_LUT4 \edb_top_inst/LUT__5071  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5071 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5072  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5072 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5073  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/n2485 ), .I3(\edb_top_inst/n2486 ), .O(\edb_top_inst/n2487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5073 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__5074  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/n2484 ), .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I3(\edb_top_inst/n2487 ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3730, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5074 .LUTMASK = 16'h3730;
    EFX_LUT4 \edb_top_inst/LUT__5075  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5075 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5076  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5076 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5077  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n20 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5077 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5078  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5078 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5079  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5079 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5080  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n10 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5080 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5081  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5081 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5082  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5082 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5083  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), .O(\edb_top_inst/n2488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5083 .LUTMASK = 16'hefef;
    EFX_LUT4 \edb_top_inst/LUT__5085  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n2490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5085 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5086  (.I0(\edb_top_inst/n2488 ), .I1(\edb_top_inst/n2490 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5086 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5087  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0909, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5087 .LUTMASK = 16'h0909;
    EFX_LUT4 \edb_top_inst/LUT__5088  (.I0(\edb_top_inst/n2490 ), .I1(\edb_top_inst/n2491 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/equal_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5088 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__5089  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5089 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__5090  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n2492 ), .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he83f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5090 .LUTMASK = 16'he83f;
    EFX_LUT4 \edb_top_inst/LUT__5091  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n2494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5091 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5092  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n2495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5092 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5093  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/n2494 ), .I3(\edb_top_inst/n2495 ), .O(\edb_top_inst/n2496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5093 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__5094  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/n2493 ), .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .I3(\edb_top_inst/n2496 ), .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3730, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5094 .LUTMASK = 16'h3730;
    EFX_LUT4 \edb_top_inst/LUT__5095  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5095 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5096  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5096 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5097  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n20 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5097 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5098  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5098 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5099  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5099 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5100  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n10 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5100 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5101  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5101 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5102  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5102 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5103  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5103 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5104  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5104 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5105  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5105 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__5106  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2497 ), .O(\edb_top_inst/n2498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5106 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__5107  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5107 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__5108  (.I0(\edb_top_inst/n2499 ), .I1(\edb_top_inst/n2498 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5108 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5109  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5109 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5110  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5110 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5111  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5111 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5112  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5112 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5113  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n2500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5113 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__5114  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n2500 ), .O(\edb_top_inst/n2501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5114 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__5115  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/n2502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5115 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__5116  (.I0(\edb_top_inst/n2502 ), .I1(\edb_top_inst/n2501 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5116 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5117  (.I0(\edb_top_inst/la0/la_trig_mask [9]), 
            .I1(\edb_top_inst/la0/la_trig_mask [10]), .I2(\edb_top_inst/la0/la_trig_mask [11]), 
            .I3(\edb_top_inst/la0/la_trig_mask [12]), .O(\edb_top_inst/n2503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5117 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5118  (.I0(\edb_top_inst/la0/la_trig_mask [0]), 
            .I1(\edb_top_inst/la0/la_trig_mask [2]), .I2(\edb_top_inst/la0/la_trig_mask [3]), 
            .I3(\edb_top_inst/la0/la_trig_mask [4]), .O(\edb_top_inst/n2504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5118 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5119  (.I0(\edb_top_inst/la0/la_trig_mask [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [6]), .I2(\edb_top_inst/n2504 ), 
            .O(\edb_top_inst/n2505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5119 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5120  (.I0(\edb_top_inst/la0/la_trig_mask [5]), 
            .I1(\edb_top_inst/la0/la_trig_mask [7]), .I2(\edb_top_inst/la0/la_trig_mask [8]), 
            .I3(\edb_top_inst/la0/la_trig_mask [13]), .O(\edb_top_inst/n2506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5120 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5121  (.I0(\edb_top_inst/la0/la_trig_mask [13]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [2]), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5121 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5122  (.I0(\edb_top_inst/la0/la_trig_mask [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [4]), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5122 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5123  (.I0(\edb_top_inst/la0/la_trig_mask [12]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [1]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5123 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5124  (.I0(\edb_top_inst/la0/la_trig_mask [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [3]), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5124 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5125  (.I0(\edb_top_inst/n2507 ), .I1(\edb_top_inst/n2508 ), 
            .I2(\edb_top_inst/n2509 ), .I3(\edb_top_inst/n2510 ), .O(\edb_top_inst/n2511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5125 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5126  (.I0(\edb_top_inst/la0/la_trig_mask [8]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [0]), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5126 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5127  (.I0(\edb_top_inst/la0/la_trig_mask [9]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [5]), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5127 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5128  (.I0(\edb_top_inst/la0/la_trig_mask [11]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [10]), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5128 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5129  (.I0(\edb_top_inst/n2511 ), .I1(\edb_top_inst/n2512 ), 
            .I2(\edb_top_inst/n2513 ), .I3(\edb_top_inst/n2514 ), .O(\edb_top_inst/n2515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5129 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5130  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [12]), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [5]), .O(\edb_top_inst/n2516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5130 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5131  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [8]), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [0]), .O(\edb_top_inst/n2517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5131 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5132  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [13]), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [4]), .O(\edb_top_inst/n2518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5132 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5133  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [6]), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [2]), .O(\edb_top_inst/n2519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5133 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5134  (.I0(\edb_top_inst/n2516 ), .I1(\edb_top_inst/n2517 ), 
            .I2(\edb_top_inst/n2518 ), .I3(\edb_top_inst/n2519 ), .O(\edb_top_inst/n2520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5134 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5135  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [10]), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [1]), .O(\edb_top_inst/n2521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5135 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5136  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [11]), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [3]), .O(\edb_top_inst/n2522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5136 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5137  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [9]), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [7]), .O(\edb_top_inst/n2523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5137 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5138  (.I0(\edb_top_inst/n2520 ), .I1(\edb_top_inst/n2521 ), 
            .I2(\edb_top_inst/n2522 ), .I3(\edb_top_inst/n2523 ), .O(\edb_top_inst/n2524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5138 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5139  (.I0(\edb_top_inst/la0/la_trig_pattern [0]), 
            .I1(\edb_top_inst/n2515 ), .I2(\edb_top_inst/n2524 ), .I3(\edb_top_inst/la0/la_trig_pattern [1]), 
            .O(\edb_top_inst/n2525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0df2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5139 .LUTMASK = 16'h0df2;
    EFX_LUT4 \edb_top_inst/LUT__5140  (.I0(\edb_top_inst/n2505 ), .I1(\edb_top_inst/n2506 ), 
            .I2(\edb_top_inst/n2503 ), .I3(\edb_top_inst/n2525 ), .O(\edb_top_inst/la0/trigger_tu/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5140 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5141  (.I0(\edb_top_inst/la0/skip_count [7]), 
            .I1(\edb_top_inst/la0/skip_count [8]), .I2(\edb_top_inst/la0/skip_count [9]), 
            .O(\edb_top_inst/n2526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5141 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5142  (.I0(\edb_top_inst/la0/skip_count [10]), 
            .I1(\edb_top_inst/la0/skip_count [11]), .I2(\edb_top_inst/la0/skip_count [12]), 
            .O(\edb_top_inst/n2527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5142 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5143  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .I2(\edb_top_inst/la0/skip_count [2]), 
            .I3(\edb_top_inst/la0/skip_count [3]), .O(\edb_top_inst/n2528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5143 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5144  (.I0(\edb_top_inst/la0/skip_count [4]), 
            .I1(\edb_top_inst/la0/skip_count [5]), .I2(\edb_top_inst/la0/skip_count [6]), 
            .O(\edb_top_inst/n2529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5144 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5145  (.I0(\edb_top_inst/n2526 ), .I1(\edb_top_inst/n2527 ), 
            .I2(\edb_top_inst/n2528 ), .I3(\edb_top_inst/n2529 ), .O(\edb_top_inst/n2530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5145 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5146  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/la0/skip_count [14]), .I2(\edb_top_inst/la0/skip_count [15]), 
            .I3(\edb_top_inst/la0/skip_count [16]), .O(\edb_top_inst/n2531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5146 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5147  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/la0/skip_count [18]), .I2(\edb_top_inst/la0/skip_count [19]), 
            .O(\edb_top_inst/n2532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5147 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5148  (.I0(\edb_top_inst/la0/skip_count [20]), 
            .I1(\edb_top_inst/la0/skip_count [21]), .I2(\edb_top_inst/n2531 ), 
            .I3(\edb_top_inst/n2532 ), .O(\edb_top_inst/n2533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5148 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5149  (.I0(\edb_top_inst/la0/skip_count [31]), 
            .I1(\edb_top_inst/la0/skip_count [32]), .I2(\edb_top_inst/la0/skip_count [33]), 
            .I3(\edb_top_inst/la0/skip_count [34]), .O(\edb_top_inst/n2534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5149 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5150  (.I0(\edb_top_inst/la0/skip_count [35]), 
            .I1(\edb_top_inst/la0/skip_count [36]), .I2(\edb_top_inst/la0/skip_count [37]), 
            .O(\edb_top_inst/n2535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5150 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5151  (.I0(\edb_top_inst/la0/skip_count [38]), 
            .I1(\edb_top_inst/la0/skip_count [39]), .I2(\edb_top_inst/n2534 ), 
            .I3(\edb_top_inst/n2535 ), .O(\edb_top_inst/n2536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5151 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5152  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/skip_count [23]), .I2(\edb_top_inst/la0/skip_count [24]), 
            .I3(\edb_top_inst/la0/skip_count [25]), .O(\edb_top_inst/n2537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5152 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5153  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/skip_count [27]), .I2(\edb_top_inst/la0/skip_count [28]), 
            .I3(\edb_top_inst/la0/skip_count [29]), .O(\edb_top_inst/n2538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5153 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5154  (.I0(\edb_top_inst/la0/skip_count [30]), 
            .I1(\edb_top_inst/n2537 ), .I2(\edb_top_inst/n2538 ), .O(\edb_top_inst/n2539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5154 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5155  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2533 ), 
            .I2(\edb_top_inst/n2536 ), .I3(\edb_top_inst/n2539 ), .O(\edb_top_inst/n2540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5155 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5156  (.I0(\edb_top_inst/la0/skip_count [41]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41]), 
            .O(\edb_top_inst/n2541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5156 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5157  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/n2541 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40]), 
            .I3(\edb_top_inst/n2540 ), .O(\edb_top_inst/n2542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5157 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5158  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2533 ), 
            .I2(\edb_top_inst/n2537 ), .O(\edb_top_inst/n2543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5158 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5159  (.I0(\edb_top_inst/la0/skip_count [27]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27]), 
            .O(\edb_top_inst/n2544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5159 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5160  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/n2544 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26]), 
            .I3(\edb_top_inst/n2543 ), .O(\edb_top_inst/n2545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5160 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5161  (.I0(\edb_top_inst/n2542 ), .I1(\edb_top_inst/n2545 ), 
            .O(\edb_top_inst/n2546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5161 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5162  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17]), 
            .O(\edb_top_inst/n2547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5162 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5163  (.I0(\edb_top_inst/la0/skip_count [18]), 
            .I1(\edb_top_inst/la0/skip_count [19]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18]), 
            .O(\edb_top_inst/n2548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5163 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5164  (.I0(\edb_top_inst/la0/skip_count [18]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18]), 
            .I2(\edb_top_inst/la0/skip_count [19]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19]), 
            .O(\edb_top_inst/n2549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5164 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5165  (.I0(\edb_top_inst/n2548 ), .I1(\edb_top_inst/n2549 ), 
            .I2(\edb_top_inst/la0/skip_count [17]), .I3(\edb_top_inst/n2547 ), 
            .O(\edb_top_inst/n2550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a33, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5165 .LUTMASK = 16'h3a33;
    EFX_LUT4 \edb_top_inst/LUT__5166  (.I0(\edb_top_inst/la0/skip_count [21]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21]), 
            .O(\edb_top_inst/n2551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5166 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5167  (.I0(\edb_top_inst/n2551 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20]), 
            .I2(\edb_top_inst/la0/skip_count [20]), .O(\edb_top_inst/n2552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5167 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5168  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2531 ), 
            .I2(\edb_top_inst/n2552 ), .I3(\edb_top_inst/n2547 ), .O(\edb_top_inst/n2553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h778f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5168 .LUTMASK = 16'h778f;
    EFX_LUT4 \edb_top_inst/LUT__5169  (.I0(\edb_top_inst/la0/skip_count [20]), 
            .I1(\edb_top_inst/n2551 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20]), 
            .I3(\edb_top_inst/n2532 ), .O(\edb_top_inst/n2554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5169 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5170  (.I0(\edb_top_inst/n2547 ), .I1(\edb_top_inst/n2554 ), 
            .I2(\edb_top_inst/n2550 ), .I3(\edb_top_inst/n2553 ), .O(\edb_top_inst/n2555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5170 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__5171  (.I0(\edb_top_inst/la0/skip_count [39]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39]), 
            .O(\edb_top_inst/n2556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5171 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5172  (.I0(\edb_top_inst/la0/skip_count [38]), 
            .I1(\edb_top_inst/n2556 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .I3(\edb_top_inst/n2535 ), .O(\edb_top_inst/n2557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5172 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5173  (.I0(\edb_top_inst/la0/skip_count [36]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36]), 
            .O(\edb_top_inst/n2558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5173 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5174  (.I0(\edb_top_inst/n2557 ), .I1(\edb_top_inst/n2558 ), 
            .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35]), 
            .I3(\edb_top_inst/la0/skip_count [35]), .O(\edb_top_inst/n2559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5174 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__5175  (.I0(\edb_top_inst/n2558 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .I2(\edb_top_inst/la0/skip_count [38]), .O(\edb_top_inst/n2560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5175 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5176  (.I0(\edb_top_inst/n2556 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35]), 
            .I2(\edb_top_inst/la0/skip_count [35]), .I3(\edb_top_inst/n2560 ), 
            .O(\edb_top_inst/n2561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5176 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__5177  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2533 ), 
            .I2(\edb_top_inst/n2539 ), .O(\edb_top_inst/n2562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5177 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5178  (.I0(\edb_top_inst/n2559 ), .I1(\edb_top_inst/n2561 ), 
            .I2(\edb_top_inst/n2534 ), .I3(\edb_top_inst/n2562 ), .O(\edb_top_inst/n2563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5178 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__5179  (.I0(\edb_top_inst/la0/skip_count [33]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33]), 
            .I2(\edb_top_inst/la0/skip_count [34]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34]), 
            .O(\edb_top_inst/n2564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5179 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5180  (.I0(\edb_top_inst/la0/skip_count [33]), 
            .I1(\edb_top_inst/la0/skip_count [34]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33]), 
            .O(\edb_top_inst/n2565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5180 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5181  (.I0(\edb_top_inst/n2565 ), .I1(\edb_top_inst/n2564 ), 
            .I2(\edb_top_inst/la0/skip_count [32]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32]), 
            .O(\edb_top_inst/n2566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5181 .LUTMASK = 16'hfa3f;
    EFX_LUT4 \edb_top_inst/LUT__5182  (.I0(\edb_top_inst/la0/skip_count [32]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32]), 
            .I2(\edb_top_inst/n2564 ), .O(\edb_top_inst/n2567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5182 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__5183  (.I0(\edb_top_inst/n2566 ), .I1(\edb_top_inst/n2567 ), 
            .I2(\edb_top_inst/la0/skip_count [31]), .I3(\edb_top_inst/n2562 ), 
            .O(\edb_top_inst/n2568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5cc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5183 .LUTMASK = 16'hc5cc;
    EFX_LUT4 \edb_top_inst/LUT__5184  (.I0(\edb_top_inst/la0/skip_count [4]), 
            .I1(\edb_top_inst/n2528 ), .O(\edb_top_inst/n2569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5184 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5185  (.I0(\edb_top_inst/la0/skip_count [6]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6]), 
            .O(\edb_top_inst/n2570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5185 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5186  (.I0(\edb_top_inst/la0/skip_count [5]), 
            .I1(\edb_top_inst/n2570 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5]), 
            .I3(\edb_top_inst/n2569 ), .O(\edb_top_inst/n2571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5186 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5187  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2533 ), 
            .O(\edb_top_inst/n2572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5187 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5188  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22]), 
            .O(\edb_top_inst/n2573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5188 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5189  (.I0(\edb_top_inst/n2571 ), .I1(\edb_top_inst/n2572 ), 
            .I2(\edb_top_inst/n2573 ), .O(\edb_top_inst/n2574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5189 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5190  (.I0(\edb_top_inst/n2555 ), .I1(\edb_top_inst/n2563 ), 
            .I2(\edb_top_inst/n2568 ), .I3(\edb_top_inst/n2574 ), .O(\edb_top_inst/n2575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5190 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5191  (.I0(\edb_top_inst/la0/skip_count [23]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .I2(\edb_top_inst/la0/skip_count [30]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30]), 
            .O(\edb_top_inst/n2576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5191 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5192  (.I0(\edb_top_inst/la0/skip_count [23]), 
            .I1(\edb_top_inst/la0/skip_count [30]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .O(\edb_top_inst/n2577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4182, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5192 .LUTMASK = 16'h4182;
    EFX_LUT4 \edb_top_inst/LUT__5193  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/n2577 ), .O(\edb_top_inst/n2578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5193 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5194  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .I1(\edb_top_inst/n2537 ), .I2(\edb_top_inst/n2538 ), .I3(\edb_top_inst/n2578 ), 
            .O(\edb_top_inst/n2579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc07f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5194 .LUTMASK = 16'hc07f;
    EFX_LUT4 \edb_top_inst/LUT__5195  (.I0(\edb_top_inst/n2579 ), .I1(\edb_top_inst/la0/skip_count [22]), 
            .I2(\edb_top_inst/n2576 ), .I3(\edb_top_inst/n2572 ), .O(\edb_top_inst/n2580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd5f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5195 .LUTMASK = 16'hd5f0;
    EFX_LUT4 \edb_top_inst/LUT__5196  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/la0/skip_count [14]), .I2(\edb_top_inst/n2530 ), 
            .O(\edb_top_inst/n2581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5196 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5197  (.I0(\edb_top_inst/la0/skip_count [16]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16]), 
            .O(\edb_top_inst/n2582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5197 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5198  (.I0(\edb_top_inst/la0/skip_count [15]), 
            .I1(\edb_top_inst/n2582 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15]), 
            .I3(\edb_top_inst/n2581 ), .O(\edb_top_inst/n2583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5198 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5199  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/skip_count [41]), .I2(\edb_top_inst/la0/skip_count [42]), 
            .I3(\edb_top_inst/la0/skip_count [43]), .O(\edb_top_inst/n2584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5199 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5200  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/la0/skip_count [45]), .I2(\edb_top_inst/la0/skip_count [46]), 
            .I3(\edb_top_inst/la0/skip_count [47]), .O(\edb_top_inst/n2585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5200 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5201  (.I0(\edb_top_inst/la0/skip_count [48]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48]), 
            .O(\edb_top_inst/n2586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5201 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5202  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2584 ), 
            .I2(\edb_top_inst/n2585 ), .I3(\edb_top_inst/n2586 ), .O(\edb_top_inst/n2587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5202 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__5203  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/skip_count [41]), .I2(\edb_top_inst/la0/skip_count [42]), 
            .O(\edb_top_inst/n2588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5203 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5204  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2588 ), 
            .I2(\edb_top_inst/la0/skip_count [43]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43]), 
            .O(\edb_top_inst/n2589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8778, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5204 .LUTMASK = 16'h8778;
    EFX_LUT4 \edb_top_inst/LUT__5205  (.I0(\edb_top_inst/n2583 ), .I1(\edb_top_inst/n2587 ), 
            .I2(\edb_top_inst/n2589 ), .I3(\edb_top_inst/n2580 ), .O(\edb_top_inst/n2590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5205 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5206  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/skip_count [27]), .I2(\edb_top_inst/n2537 ), 
            .O(\edb_top_inst/n2591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5206 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5207  (.I0(\edb_top_inst/n2530 ), .I1(\edb_top_inst/n2533 ), 
            .I2(\edb_top_inst/n2591 ), .O(\edb_top_inst/n2592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5207 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5208  (.I0(\edb_top_inst/la0/skip_count [29]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29]), 
            .O(\edb_top_inst/n2593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5208 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5209  (.I0(\edb_top_inst/la0/skip_count [28]), 
            .I1(\edb_top_inst/n2593 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28]), 
            .I3(\edb_top_inst/n2592 ), .O(\edb_top_inst/n2594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5209 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5210  (.I0(\edb_top_inst/la0/skip_count [47]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47]), 
            .O(\edb_top_inst/n2595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5210 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5211  (.I0(\edb_top_inst/la0/skip_count [46]), 
            .I1(\edb_top_inst/la0/skip_count [45]), .I2(\edb_top_inst/n2595 ), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45]), 
            .O(\edb_top_inst/n2596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5211 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__5212  (.I0(\edb_top_inst/n2595 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45]), 
            .I2(\edb_top_inst/la0/skip_count [45]), .O(\edb_top_inst/n2597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5212 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5213  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/n2584 ), .O(\edb_top_inst/n2598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5213 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5214  (.I0(\edb_top_inst/n2596 ), .I1(\edb_top_inst/n2597 ), 
            .I2(\edb_top_inst/n2540 ), .I3(\edb_top_inst/n2598 ), .O(\edb_top_inst/n2599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5214 .LUTMASK = 16'h5ccc;
    EFX_LUT4 \edb_top_inst/LUT__5215  (.I0(\edb_top_inst/n2526 ), .I1(\edb_top_inst/n2528 ), 
            .I2(\edb_top_inst/n2529 ), .O(\edb_top_inst/n2600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5215 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5216  (.I0(\edb_top_inst/la0/skip_count [10]), 
            .I1(\edb_top_inst/n2600 ), .O(\edb_top_inst/n2601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5216 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5217  (.I0(\edb_top_inst/la0/skip_count [12]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12]), 
            .O(\edb_top_inst/n2602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5217 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5218  (.I0(\edb_top_inst/la0/skip_count [11]), 
            .I1(\edb_top_inst/n2602 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11]), 
            .I3(\edb_top_inst/n2601 ), .O(\edb_top_inst/n2603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5218 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5219  (.I0(\edb_top_inst/la0/skip_count [14]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14]), 
            .O(\edb_top_inst/n2604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5219 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5220  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/n2604 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13]), 
            .I3(\edb_top_inst/n2530 ), .O(\edb_top_inst/n2605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5220 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5221  (.I0(\edb_top_inst/la0/skip_count [7]), 
            .I1(\edb_top_inst/n2528 ), .I2(\edb_top_inst/n2529 ), .O(\edb_top_inst/n2606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5221 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5222  (.I0(\edb_top_inst/la0/skip_count [9]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9]), 
            .O(\edb_top_inst/n2607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5222 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5223  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/n2607 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8]), 
            .I3(\edb_top_inst/n2606 ), .O(\edb_top_inst/n2608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5223 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5224  (.I0(\edb_top_inst/n2528 ), .I1(\edb_top_inst/n2529 ), 
            .O(\edb_top_inst/n2609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5224 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5225  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .O(\edb_top_inst/n2610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5225 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5226  (.I0(\edb_top_inst/n2610 ), .I1(\edb_top_inst/la0/skip_count [4]), 
            .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4]), 
            .I3(\edb_top_inst/n2528 ), .O(\edb_top_inst/n2611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5226 .LUTMASK = 16'h1441;
    EFX_LUT4 \edb_top_inst/LUT__5227  (.I0(\edb_top_inst/la0/skip_count [7]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7]), 
            .I2(\edb_top_inst/n2609 ), .I3(\edb_top_inst/n2611 ), .O(\edb_top_inst/n2612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5227 .LUTMASK = 16'h6900;
    EFX_LUT4 \edb_top_inst/LUT__5228  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .O(\edb_top_inst/n2613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5228 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5229  (.I0(\edb_top_inst/la0/skip_count [3]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3]), 
            .O(\edb_top_inst/n2614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5229 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5230  (.I0(\edb_top_inst/la0/skip_count [2]), 
            .I1(\edb_top_inst/n2614 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2]), 
            .I3(\edb_top_inst/n2613 ), .O(\edb_top_inst/n2615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5230 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5231  (.I0(\edb_top_inst/n2615 ), .I1(\edb_top_inst/la0/skip_count [10]), 
            .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10]), 
            .I3(\edb_top_inst/n2600 ), .O(\edb_top_inst/n2616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5231 .LUTMASK = 16'h1441;
    EFX_LUT4 \edb_top_inst/LUT__5232  (.I0(\edb_top_inst/n2605 ), .I1(\edb_top_inst/n2608 ), 
            .I2(\edb_top_inst/n2612 ), .I3(\edb_top_inst/n2616 ), .O(\edb_top_inst/n2617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5232 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5233  (.I0(\edb_top_inst/n2594 ), .I1(\edb_top_inst/n2603 ), 
            .I2(\edb_top_inst/n2599 ), .I3(\edb_top_inst/n2617 ), .O(\edb_top_inst/n2618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5233 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5234  (.I0(\edb_top_inst/n2546 ), .I1(\edb_top_inst/n2575 ), 
            .I2(\edb_top_inst/n2590 ), .I3(\edb_top_inst/n2618 ), .O(\edb_top_inst/n2619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5234 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5235  (.I0(\edb_top_inst/la0/skip_count [48]), 
            .I1(\edb_top_inst/n2584 ), .I2(\edb_top_inst/n2585 ), .O(\edb_top_inst/n2620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5235 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5236  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/n2540 ), .I2(\edb_top_inst/n2620 ), .O(\edb_top_inst/n2621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5236 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5237  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/skip_count [50]), .I2(\edb_top_inst/la0/skip_count [51]), 
            .O(\edb_top_inst/n2622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5237 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5238  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52]), 
            .O(\edb_top_inst/n2623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5238 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5239  (.I0(\edb_top_inst/la0/skip_count [50]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50]), 
            .O(\edb_top_inst/n2624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5239 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5240  (.I0(\edb_top_inst/n2622 ), .I1(\edb_top_inst/n2623 ), 
            .I2(\edb_top_inst/n2621 ), .I3(\edb_top_inst/n2624 ), .O(\edb_top_inst/n2625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5240 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__5241  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/la0/skip_count [53]), .I2(\edb_top_inst/la0/skip_count [54]), 
            .I3(\edb_top_inst/n2622 ), .O(\edb_top_inst/n2626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5241 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5242  (.I0(\edb_top_inst/n2620 ), .I1(\edb_top_inst/n2626 ), 
            .O(\edb_top_inst/n2627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5242 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5243  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2627 ), 
            .I2(\edb_top_inst/la0/skip_count [55]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55]), 
            .O(\edb_top_inst/n2628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8778, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5243 .LUTMASK = 16'h8778;
    EFX_LUT4 \edb_top_inst/LUT__5244  (.I0(\edb_top_inst/la0/skip_count [35]), 
            .I1(\edb_top_inst/la0/skip_count [36]), .I2(\edb_top_inst/n2534 ), 
            .O(\edb_top_inst/n2629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5244 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5245  (.I0(\edb_top_inst/la0/skip_count [31]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31]), 
            .O(\edb_top_inst/n2630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5245 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5246  (.I0(\edb_top_inst/la0/skip_count [37]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37]), 
            .O(\edb_top_inst/n2631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5246 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5247  (.I0(\edb_top_inst/n2629 ), .I1(\edb_top_inst/n2631 ), 
            .I2(\edb_top_inst/n2630 ), .I3(\edb_top_inst/n2562 ), .O(\edb_top_inst/n2632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5247 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__5248  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58]), 
            .O(\edb_top_inst/n2633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5248 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5249  (.I0(\edb_top_inst/la0/skip_count [57]), 
            .I1(\edb_top_inst/la0/skip_count [56]), .I2(\edb_top_inst/n2633 ), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .O(\edb_top_inst/n2634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5249 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__5250  (.I0(\edb_top_inst/n2633 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .I2(\edb_top_inst/la0/skip_count [56]), .O(\edb_top_inst/n2635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5250 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5251  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/n2620 ), .I2(\edb_top_inst/n2626 ), .O(\edb_top_inst/n2636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5251 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5252  (.I0(\edb_top_inst/n2634 ), .I1(\edb_top_inst/n2635 ), 
            .I2(\edb_top_inst/n2540 ), .I3(\edb_top_inst/n2636 ), .O(\edb_top_inst/n2637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5252 .LUTMASK = 16'h5ccc;
    EFX_LUT4 \edb_top_inst/LUT__5253  (.I0(\edb_top_inst/n2628 ), .I1(\edb_top_inst/n2632 ), 
            .I2(\edb_top_inst/n2637 ), .O(\edb_top_inst/n2638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5253 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5254  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/skip_count [23]), .I2(\edb_top_inst/n2530 ), 
            .I3(\edb_top_inst/n2533 ), .O(\edb_top_inst/n2639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5254 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5255  (.I0(\edb_top_inst/la0/skip_count [25]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25]), 
            .O(\edb_top_inst/n2640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5255 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5256  (.I0(\edb_top_inst/la0/skip_count [24]), 
            .I1(\edb_top_inst/n2640 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24]), 
            .I3(\edb_top_inst/n2639 ), .O(\edb_top_inst/n2641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5256 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5257  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/la0/skip_count [56]), .O(\edb_top_inst/n2642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5257 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5258  (.I0(\edb_top_inst/la0/skip_count [57]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57]), 
            .O(\edb_top_inst/n2643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5258 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5259  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2627 ), 
            .I2(\edb_top_inst/n2642 ), .I3(\edb_top_inst/n2643 ), .O(\edb_top_inst/n2644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5259 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__5260  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/la0/skip_count [56]), .I2(\edb_top_inst/la0/skip_count [57]), 
            .I3(\edb_top_inst/la0/skip_count [58]), .O(\edb_top_inst/n2645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5260 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5261  (.I0(\edb_top_inst/la0/skip_count [59]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59]), 
            .O(\edb_top_inst/n2646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5261 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5262  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2627 ), 
            .I2(\edb_top_inst/n2645 ), .I3(\edb_top_inst/n2646 ), .O(\edb_top_inst/n2647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5262 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__5263  (.I0(\edb_top_inst/la0/skip_count [59]), 
            .I1(\edb_top_inst/n2620 ), .I2(\edb_top_inst/n2626 ), .I3(\edb_top_inst/n2645 ), 
            .O(\edb_top_inst/n2648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5263 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5264  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2648 ), 
            .I2(\edb_top_inst/la0/skip_count [60]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60]), 
            .O(\edb_top_inst/n2649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8778, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5264 .LUTMASK = 16'h8778;
    EFX_LUT4 \edb_top_inst/LUT__5265  (.I0(\edb_top_inst/n2641 ), .I1(\edb_top_inst/n2644 ), 
            .I2(\edb_top_inst/n2647 ), .I3(\edb_top_inst/n2649 ), .O(\edb_top_inst/n2650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5265 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5266  (.I0(\edb_top_inst/la0/skip_count [59]), 
            .I1(\edb_top_inst/la0/skip_count [60]), .I2(\edb_top_inst/n2645 ), 
            .O(\edb_top_inst/n2651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5266 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5267  (.I0(\edb_top_inst/la0/skip_count [61]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61]), 
            .O(\edb_top_inst/n2652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5267 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5268  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/skip_count [50]), .O(\edb_top_inst/n2653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5268 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5269  (.I0(\edb_top_inst/la0/skip_count [51]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .I2(\edb_top_inst/n2653 ), .O(\edb_top_inst/n2654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5269 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__5270  (.I0(\edb_top_inst/n2626 ), .I1(\edb_top_inst/n2651 ), 
            .I2(\edb_top_inst/n2652 ), .I3(\edb_top_inst/n2654 ), .O(\edb_top_inst/n2655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5270 .LUTMASK = 16'h8700;
    EFX_LUT4 \edb_top_inst/LUT__5271  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2620 ), 
            .I2(\edb_top_inst/n2655 ), .O(\edb_top_inst/n2656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5271 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5272  (.I0(\edb_top_inst/n2652 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .I2(\edb_top_inst/la0/skip_count [51]), .O(\edb_top_inst/n2657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5272 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5273  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2620 ), 
            .I2(\edb_top_inst/n2653 ), .I3(\edb_top_inst/n2657 ), .O(\edb_top_inst/n2658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5273 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5274  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49]), 
            .O(\edb_top_inst/n2659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5274 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5275  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .I2(\edb_top_inst/la0/skip_count [46]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .O(\edb_top_inst/n2660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5275 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5276  (.I0(\edb_top_inst/n2659 ), .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42]), 
            .I2(\edb_top_inst/la0/skip_count [42]), .I3(\edb_top_inst/n2660 ), 
            .O(\edb_top_inst/n2661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5276 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__5277  (.I0(\edb_top_inst/la0/skip_count [41]), 
            .I1(\edb_top_inst/la0/skip_count [40]), .I2(\edb_top_inst/n2540 ), 
            .I3(\edb_top_inst/n2661 ), .O(\edb_top_inst/n2662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5277 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__5278  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .I1(\edb_top_inst/la0/skip_count [46]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .I3(\edb_top_inst/la0/skip_count [44]), .O(\edb_top_inst/n2663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5278 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__5279  (.I0(\edb_top_inst/la0/skip_count [45]), 
            .I1(\edb_top_inst/la0/skip_count [46]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .O(\edb_top_inst/n2664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5279 .LUTMASK = 16'h9696;
    EFX_LUT4 \edb_top_inst/LUT__5280  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/n2664 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .O(\edb_top_inst/n2665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5280 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5281  (.I0(\edb_top_inst/n2665 ), .I1(\edb_top_inst/n2663 ), 
            .I2(\edb_top_inst/n2660 ), .I3(\edb_top_inst/n2584 ), .O(\edb_top_inst/n2666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5281 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__5282  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/skip_count [41]), .I2(\edb_top_inst/la0/skip_count [42]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42]), 
            .O(\edb_top_inst/n2667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5282 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__5283  (.I0(\edb_top_inst/n2620 ), .I1(\edb_top_inst/n2659 ), 
            .I2(\edb_top_inst/n2667 ), .O(\edb_top_inst/n2668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5283 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__5284  (.I0(\edb_top_inst/n2540 ), .I1(\edb_top_inst/n2666 ), 
            .I2(\edb_top_inst/n2668 ), .O(\edb_top_inst/n2669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5284 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5285  (.I0(\edb_top_inst/n2662 ), .I1(\edb_top_inst/n2669 ), 
            .I2(\edb_top_inst/n2656 ), .I3(\edb_top_inst/n2658 ), .O(\edb_top_inst/n2670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5285 .LUTMASK = 16'heee0;
    EFX_LUT4 \edb_top_inst/LUT__5286  (.I0(\edb_top_inst/n2625 ), .I1(\edb_top_inst/n2638 ), 
            .I2(\edb_top_inst/n2650 ), .I3(\edb_top_inst/n2670 ), .O(\edb_top_inst/n2671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5286 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5287  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/n2540 ), .I2(\edb_top_inst/n2620 ), .I3(\edb_top_inst/n2622 ), 
            .O(\edb_top_inst/n2672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5287 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5288  (.I0(\edb_top_inst/la0/skip_count [54]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54]), 
            .O(\edb_top_inst/n2673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5288 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5289  (.I0(\edb_top_inst/la0/skip_count [53]), 
            .I1(\edb_top_inst/n2673 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53]), 
            .I3(\edb_top_inst/n2672 ), .O(\edb_top_inst/n2674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5289 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5290  (.I0(\edb_top_inst/la0/skip_count [61]), 
            .I1(\edb_top_inst/n2540 ), .I2(\edb_top_inst/n2627 ), .I3(\edb_top_inst/n2651 ), 
            .O(\edb_top_inst/n2675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5290 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5291  (.I0(\edb_top_inst/la0/skip_count [63]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63]), 
            .O(\edb_top_inst/n2676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5291 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5292  (.I0(\edb_top_inst/la0/skip_count [62]), 
            .I1(\edb_top_inst/n2676 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62]), 
            .I3(\edb_top_inst/n2675 ), .O(\edb_top_inst/n2677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5292 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5293  (.I0(\edb_top_inst/n2674 ), .I1(\edb_top_inst/n2677 ), 
            .O(\edb_top_inst/n2678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5293 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5294  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5294 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__5295  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/n2678 ), .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/n2671 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5295 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5296  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [1]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5296 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5297  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [2]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5297 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5298  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [3]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5298 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5299  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [4]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5299 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5300  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [5]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5300 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5301  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [6]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5301 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5302  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [7]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5302 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5303  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [8]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5303 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5304  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [9]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5304 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5305  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [10]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5305 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5306  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [11]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5306 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5307  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [12]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5307 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5308  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [13]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5308 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5309  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [14]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5309 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5310  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [15]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5310 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5311  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [16]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5311 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5312  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [17]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5312 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5313  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [18]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5313 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5314  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [19]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5314 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5315  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [20]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5315 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5316  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [21]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5316 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5317  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [22]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5317 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5318  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [23]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5318 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5319  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [24]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5319 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5320  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [25]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5320 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5321  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [26]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5321 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5322  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [27]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5322 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5323  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [28]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5323 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5324  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [29]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5324 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5325  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [30]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5325 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5326  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [31]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5326 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5327  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [32]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5327 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5328  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [33]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5328 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5329  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [34]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5329 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5330  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [35]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5330 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5331  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [36]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5331 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5332  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [37]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5332 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5333  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [38]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5333 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5334  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [39]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5334 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5335  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [40]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5335 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5336  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [41]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5336 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5337  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [42]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5337 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5338  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [43]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5338 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5339  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [44]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5339 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5340  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [45]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5340 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5341  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [46]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5341 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5342  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [47]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5342 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5343  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [48]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5343 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5344  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [49]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5344 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5345  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [50]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5345 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5346  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [51]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5346 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5347  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [52]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5347 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5348  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [53]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5348 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5349  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [54]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5349 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5350  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [55]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5350 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5351  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [56]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5351 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5352  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [57]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5352 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5353  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [58]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5353 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5354  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [59]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5354 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5355  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [60]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5355 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5356  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [61]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5356 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5357  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [62]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5357 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5358  (.I0(\edb_top_inst/n2671 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/trigger_skipper_n/n73 [63]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5358 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5359  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5359 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5360  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(\edb_top_inst/n2679 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .O(\edb_top_inst/n2680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5360 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__5361  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n2681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5361 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5362  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/n2681 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .O(\edb_top_inst/n2682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d82, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5362 .LUTMASK = 16'h7d82;
    EFX_LUT4 \edb_top_inst/LUT__5363  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .O(\edb_top_inst/n2683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5363 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5364  (.I0(\edb_top_inst/n2682 ), .I1(\edb_top_inst/n2680 ), 
            .I2(\edb_top_inst/n2683 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .O(\edb_top_inst/n2684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h31cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5364 .LUTMASK = 16'h31cf;
    EFX_LUT4 \edb_top_inst/LUT__5365  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n2685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5365 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5366  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .I2(\edb_top_inst/n2679 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .O(\edb_top_inst/n2686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5366 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__5367  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5367 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__5368  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/n2683 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), .O(\edb_top_inst/n2688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0df2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5368 .LUTMASK = 16'h0df2;
    EFX_LUT4 \edb_top_inst/LUT__5369  (.I0(\edb_top_inst/n2688 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/n2687 ), .I3(\edb_top_inst/n2686 ), .O(\edb_top_inst/n2689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5369 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__5370  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/n2679 ), .O(\edb_top_inst/n2690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5370 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__5371  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5371 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__5372  (.I0(\edb_top_inst/n2690 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), 
            .I2(\edb_top_inst/n2691 ), .O(\edb_top_inst/n2692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5372 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__5373  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .O(\edb_top_inst/n2693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5373 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5374  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/n2693 ), 
            .O(\edb_top_inst/n2694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5374 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5375  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .O(\edb_top_inst/n2695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5375 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5376  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I1(\edb_top_inst/n2695 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
            .O(\edb_top_inst/n2696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5376 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__5377  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n2697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5377 .LUTMASK = 16'hfe00;
    EFX_LUT4 \edb_top_inst/LUT__5378  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/n2697 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .O(\edb_top_inst/n2698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1e1e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5378 .LUTMASK = 16'h1e1e;
    EFX_LUT4 \edb_top_inst/LUT__5379  (.I0(\edb_top_inst/n2696 ), .I1(\edb_top_inst/n2698 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), .I3(\edb_top_inst/n2694 ), 
            .O(\edb_top_inst/n2699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5379 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__5380  (.I0(\edb_top_inst/n2684 ), .I1(\edb_top_inst/n2689 ), 
            .I2(\edb_top_inst/n2692 ), .I3(\edb_top_inst/n2699 ), .O(\edb_top_inst/n2700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5380 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5381  (.I0(\edb_top_inst/n2681 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/n2679 ), .I3(\edb_top_inst/la0/la_trig_pos [4]), 
            .O(\edb_top_inst/n2701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb06f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5381 .LUTMASK = 16'hb06f;
    EFX_LUT4 \edb_top_inst/LUT__5382  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .I3(\edb_top_inst/n2681 ), .O(\edb_top_inst/n2702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5415, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5382 .LUTMASK = 16'h5415;
    EFX_LUT4 \edb_top_inst/LUT__5383  (.I0(\edb_top_inst/n2701 ), .I1(\edb_top_inst/la0/la_trig_pos [12]), 
            .I2(\edb_top_inst/n2702 ), .O(\edb_top_inst/n2703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5383 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__5384  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .I2(\edb_top_inst/n2679 ), .I3(\edb_top_inst/la0/la_trig_pos [6]), 
            .O(\edb_top_inst/n2704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5384 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__5385  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n2705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5385 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5386  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/n2705 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_trig_pos [13]), .O(\edb_top_inst/n2706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5386 .LUTMASK = 16'h07f8;
    EFX_LUT4 \edb_top_inst/LUT__5387  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5387 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5388  (.I0(\edb_top_inst/la0/la_trig_pos [1]), 
            .I1(\edb_top_inst/la0/la_trig_pos [5]), .I2(\edb_top_inst/n2691 ), 
            .I3(\edb_top_inst/n2707 ), .O(\edb_top_inst/n2708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5388 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__5389  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_trig_pos [7]), .I2(\edb_top_inst/n2679 ), 
            .O(\edb_top_inst/n2709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5389 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__5390  (.I0(\edb_top_inst/n2706 ), .I1(\edb_top_inst/n2704 ), 
            .I2(\edb_top_inst/n2708 ), .I3(\edb_top_inst/n2709 ), .O(\edb_top_inst/n2710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5390 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5391  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/n2693 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [2]), .O(\edb_top_inst/n2711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5391 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__5392  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5392 .LUTMASK = 16'hfe00;
    EFX_LUT4 \edb_top_inst/LUT__5393  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_trig_pos [11]), .O(\edb_top_inst/n2713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5393 .LUTMASK = 16'h07f8;
    EFX_LUT4 \edb_top_inst/LUT__5394  (.I0(\edb_top_inst/n2712 ), .I1(\edb_top_inst/n2713 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [3]), .I3(\edb_top_inst/n2693 ), 
            .O(\edb_top_inst/n2714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5394 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__5395  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/n2705 ), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/la0/la_trig_pos [14]), 
            .O(\edb_top_inst/n2715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5395 .LUTMASK = 16'h07f8;
    EFX_LUT4 \edb_top_inst/LUT__5396  (.I0(\edb_top_inst/n2715 ), .I1(\edb_top_inst/n2714 ), 
            .I2(\edb_top_inst/n2711 ), .O(\edb_top_inst/n2716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5396 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5397  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/n2683 ), .O(\edb_top_inst/n2717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5397 .LUTMASK = 16'h0e03;
    EFX_LUT4 \edb_top_inst/LUT__5398  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [4]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5398 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5399  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/n2718 ), 
            .I3(\edb_top_inst/la0/la_trig_pos [10]), .O(\edb_top_inst/n2719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5399 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__5400  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_trig_pos [16]), .I2(\edb_top_inst/la0/la_trig_pos [15]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n2720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5400 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__5401  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/n2697 ), .I2(\edb_top_inst/n2720 ), .I3(\edb_top_inst/la0/la_trig_pos [8]), 
            .O(\edb_top_inst/n2721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5401 .LUTMASK = 16'h0e01;
    EFX_LUT4 \edb_top_inst/LUT__5402  (.I0(\edb_top_inst/la0/la_trig_pos [9]), 
            .I1(\edb_top_inst/n2719 ), .I2(\edb_top_inst/n2717 ), .I3(\edb_top_inst/n2721 ), 
            .O(\edb_top_inst/n2722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5402 .LUTMASK = 16'h1800;
    EFX_LUT4 \edb_top_inst/LUT__5403  (.I0(\edb_top_inst/n2703 ), .I1(\edb_top_inst/n2710 ), 
            .I2(\edb_top_inst/n2716 ), .I3(\edb_top_inst/n2722 ), .O(\edb_top_inst/n2723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5403 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5404  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), .O(\edb_top_inst/n2724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3fd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5404 .LUTMASK = 16'he3fd;
    EFX_LUT4 \edb_top_inst/LUT__5405  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), .I2(\edb_top_inst/n2724 ), 
            .I3(\edb_top_inst/n2693 ), .O(\edb_top_inst/n2725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5405 .LUTMASK = 16'hf077;
    EFX_LUT4 \edb_top_inst/LUT__5406  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/n2695 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), .O(\edb_top_inst/n2726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h41be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5406 .LUTMASK = 16'h41be;
    EFX_LUT4 \edb_top_inst/LUT__5407  (.I0(\edb_top_inst/n2695 ), .I1(\edb_top_inst/n2679 ), 
            .I2(\edb_top_inst/n2726 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .O(\edb_top_inst/n2727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5407 .LUTMASK = 16'h0b04;
    EFX_LUT4 \edb_top_inst/LUT__5408  (.I0(\edb_top_inst/n2695 ), .I1(\edb_top_inst/n2691 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), .O(\edb_top_inst/n2728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5408 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__5409  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/la0/la_window_depth [1]), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [0]), 
            .O(\edb_top_inst/n2729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2aa8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5409 .LUTMASK = 16'h2aa8;
    EFX_LUT4 \edb_top_inst/LUT__5410  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .I1(\edb_top_inst/n2729 ), .I2(\edb_top_inst/n2682 ), .O(\edb_top_inst/n2730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5410 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__5411  (.I0(\edb_top_inst/n2725 ), .I1(\edb_top_inst/n2728 ), 
            .I2(\edb_top_inst/n2727 ), .I3(\edb_top_inst/n2730 ), .O(\edb_top_inst/n2731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5411 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5412  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/n2718 ), 
            .O(\edb_top_inst/n2732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5412 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5413  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/n2732 ), .I3(\edb_top_inst/n2717 ), .O(\edb_top_inst/n2733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5413 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__5414  (.I0(\edb_top_inst/n2681 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), .I3(\edb_top_inst/n2694 ), 
            .O(\edb_top_inst/n2734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5414 .LUTMASK = 16'h7ecf;
    EFX_LUT4 \edb_top_inst/LUT__5415  (.I0(\edb_top_inst/n2733 ), .I1(\edb_top_inst/n2734 ), 
            .O(\edb_top_inst/n2735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5415 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5416  (.I0(\edb_top_inst/n2731 ), .I1(\edb_top_inst/n2735 ), 
            .I2(\edb_top_inst/n2700 ), .I3(\edb_top_inst/n2723 ), .O(\edb_top_inst/n2736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5416 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__5417  (.I0(\edb_top_inst/la0/la_trig_pos [11]), 
            .I1(\edb_top_inst/la0/la_trig_pos [12]), .I2(\edb_top_inst/la0/la_trig_pos [15]), 
            .I3(\edb_top_inst/la0/la_trig_pos [16]), .O(\edb_top_inst/n2737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5417 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5418  (.I0(\edb_top_inst/la0/la_trig_pos [10]), 
            .I1(\edb_top_inst/la0/la_trig_pos [13]), .I2(\edb_top_inst/la0/la_trig_pos [14]), 
            .I3(\edb_top_inst/n2737 ), .O(\edb_top_inst/n2738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5418 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5419  (.I0(\edb_top_inst/la0/la_trig_pos [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [4]), .I2(\edb_top_inst/la0/la_trig_pos [5]), 
            .I3(\edb_top_inst/la0/la_trig_pos [6]), .O(\edb_top_inst/n2739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5419 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5420  (.I0(\edb_top_inst/la0/la_trig_pos [3]), 
            .I1(\edb_top_inst/la0/la_trig_pos [7]), .I2(\edb_top_inst/la0/la_trig_pos [8]), 
            .I3(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n2740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5420 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5421  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_trig_pos [1]), .I2(\edb_top_inst/n2740 ), 
            .O(\edb_top_inst/n2741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5421 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5422  (.I0(\edb_top_inst/n2738 ), .I1(\edb_top_inst/n2739 ), 
            .I2(\edb_top_inst/n2741 ), .O(\edb_top_inst/n2742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5422 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5423  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .I2(\edb_top_inst/la0/la_num_trigger [2]), 
            .I3(\edb_top_inst/la0/la_num_trigger [3]), .O(\edb_top_inst/n2743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5423 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5424  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/n2743 ), .O(\edb_top_inst/n2744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5424 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5425  (.I0(\edb_top_inst/la0/la_num_trigger [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), .O(\edb_top_inst/n2745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5425 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5426  (.I0(\edb_top_inst/la0/la_num_trigger [5]), 
            .I1(\edb_top_inst/n2745 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I3(\edb_top_inst/n2744 ), .O(\edb_top_inst/n2746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5426 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5427  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/la0/la_num_trigger [5]), .I2(\edb_top_inst/la0/la_num_trigger [6]), 
            .O(\edb_top_inst/n2747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5427 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5428  (.I0(\edb_top_inst/la0/la_num_trigger [7]), 
            .I1(\edb_top_inst/la0/la_num_trigger [8]), .I2(\edb_top_inst/n2743 ), 
            .I3(\edb_top_inst/n2747 ), .O(\edb_top_inst/n2748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5428 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5429  (.I0(\edb_top_inst/la0/la_num_trigger [9]), 
            .I1(\edb_top_inst/la0/la_num_trigger [10]), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I3(\edb_top_inst/n2748 ), .O(\edb_top_inst/n2749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5429 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5430  (.I0(\edb_top_inst/n2743 ), .I1(\edb_top_inst/n2747 ), 
            .O(\edb_top_inst/n2750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5430 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5431  (.I0(\edb_top_inst/la0/la_num_trigger [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), .O(\edb_top_inst/n2751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5431 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5432  (.I0(\edb_top_inst/la0/la_num_trigger [7]), 
            .I1(\edb_top_inst/n2751 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I3(\edb_top_inst/n2750 ), .O(\edb_top_inst/n2752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5432 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5433  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .O(\edb_top_inst/n2753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5433 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5434  (.I0(\edb_top_inst/la0/la_num_trigger [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), .O(\edb_top_inst/n2754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5434 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5435  (.I0(\edb_top_inst/la0/la_num_trigger [2]), 
            .I1(\edb_top_inst/n2754 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I3(\edb_top_inst/n2753 ), .O(\edb_top_inst/n2755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5435 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5436  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .O(\edb_top_inst/n2756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5436 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5437  (.I0(\edb_top_inst/la0/la_num_trigger [13]), 
            .I1(\edb_top_inst/la0/la_num_trigger [14]), .I2(\edb_top_inst/la0/la_num_trigger [15]), 
            .I3(\edb_top_inst/la0/la_num_trigger [16]), .O(\edb_top_inst/n2757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5437 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5438  (.I0(\edb_top_inst/la0/la_num_trigger [11]), 
            .I1(\edb_top_inst/la0/la_num_trigger [12]), .I2(\edb_top_inst/n2757 ), 
            .O(\edb_top_inst/n2758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5438 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5439  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), .I2(\edb_top_inst/n2743 ), 
            .O(\edb_top_inst/n2759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5439 .LUTMASK = 16'h9696;
    EFX_LUT4 \edb_top_inst/LUT__5440  (.I0(\edb_top_inst/n2755 ), .I1(\edb_top_inst/n2756 ), 
            .I2(\edb_top_inst/n2759 ), .I3(\edb_top_inst/n2758 ), .O(\edb_top_inst/n2760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5440 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5441  (.I0(\edb_top_inst/n2746 ), .I1(\edb_top_inst/n2749 ), 
            .I2(\edb_top_inst/n2752 ), .I3(\edb_top_inst/n2760 ), .O(\edb_top_inst/n2761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5441 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5442  (.I0(\edb_top_inst/n2742 ), .I1(\edb_top_inst/n2761 ), 
            .O(\edb_top_inst/n2762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5442 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5443  (.I0(\edb_top_inst/la0/ts_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n2763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5443 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5444  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_trig_pos [10]), .O(\edb_top_inst/n2764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1003, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5444 .LUTMASK = 16'h1003;
    EFX_LUT4 \edb_top_inst/LUT__5445  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [4]), .I2(\edb_top_inst/la0/la_trig_pos [10]), 
            .I3(\edb_top_inst/n2764 ), .O(\edb_top_inst/n2765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5445 .LUTMASK = 16'h00fe;
    EFX_LUT4 \edb_top_inst/LUT__5446  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .I2(\edb_top_inst/la0/la_trig_pos [10]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5446 .LUTMASK = 16'h1ff0;
    EFX_LUT4 \edb_top_inst/LUT__5447  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/n2766 ), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .I3(\edb_top_inst/n2765 ), .O(\edb_top_inst/n2767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5447 .LUTMASK = 16'heee0;
    EFX_LUT4 \edb_top_inst/LUT__5448  (.I0(\edb_top_inst/la0/la_trig_pos [11]), 
            .I1(\edb_top_inst/n2681 ), .I2(\edb_top_inst/la0/la_trig_pos [12]), 
            .I3(\edb_top_inst/n2705 ), .O(\edb_top_inst/n2768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5448 .LUTMASK = 16'h7d50;
    EFX_LUT4 \edb_top_inst/LUT__5449  (.I0(\edb_top_inst/n2768 ), .I1(\edb_top_inst/la0/la_trig_pos [12]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/la0/la_trig_pos [11]), 
            .O(\edb_top_inst/n2769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h15fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5449 .LUTMASK = 16'h15fe;
    EFX_LUT4 \edb_top_inst/LUT__5450  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [7]), .I2(\edb_top_inst/la0/la_trig_pos [3]), 
            .I3(\edb_top_inst/n2679 ), .O(\edb_top_inst/n2770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5450 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__5451  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/n2683 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n2771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0df2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5451 .LUTMASK = 16'h0df2;
    EFX_LUT4 \edb_top_inst/LUT__5452  (.I0(\edb_top_inst/n2770 ), .I1(\edb_top_inst/n2771 ), 
            .I2(\edb_top_inst/n2711 ), .O(\edb_top_inst/n2772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5452 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5453  (.I0(\edb_top_inst/n2767 ), .I1(\edb_top_inst/n2769 ), 
            .I2(\edb_top_inst/n2772 ), .I3(\edb_top_inst/n2708 ), .O(\edb_top_inst/n2773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5453 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5454  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_trig_pos [14]), 
            .I3(\edb_top_inst/la0/la_trig_pos [6]), .O(\edb_top_inst/n2774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5454 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__5455  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .O(\edb_top_inst/n2775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5455 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5456  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/la0/la_trig_pos [14]), 
            .I2(\edb_top_inst/n2774 ), .O(\edb_top_inst/n2776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5456 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__5457  (.I0(\edb_top_inst/la0/la_trig_pos [14]), 
            .I1(\edb_top_inst/la0/la_trig_pos [6]), .I2(\edb_top_inst/n2775 ), 
            .I3(\edb_top_inst/n2679 ), .O(\edb_top_inst/n2777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5457 .LUTMASK = 16'hbe7f;
    EFX_LUT4 \edb_top_inst/LUT__5458  (.I0(\edb_top_inst/la0/la_trig_pos [4]), 
            .I1(\edb_top_inst/n2679 ), .O(\edb_top_inst/n2778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5458 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5459  (.I0(\edb_top_inst/n2681 ), .I1(\edb_top_inst/n2778 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [0]), .I3(\edb_top_inst/n2701 ), 
            .O(\edb_top_inst/n2779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf70f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5459 .LUTMASK = 16'hf70f;
    EFX_LUT4 \edb_top_inst/LUT__5460  (.I0(\edb_top_inst/n2706 ), .I1(\edb_top_inst/n2721 ), 
            .O(\edb_top_inst/n2780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5460 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5461  (.I0(\edb_top_inst/n2777 ), .I1(\edb_top_inst/n2776 ), 
            .I2(\edb_top_inst/n2779 ), .I3(\edb_top_inst/n2780 ), .O(\edb_top_inst/n2781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5461 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__5462  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .O(\edb_top_inst/n2782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5462 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__5463  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/n2781 ), 
            .I2(\edb_top_inst/n2773 ), .I3(\edb_top_inst/n2782 ), .O(\edb_top_inst/n2783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5463 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__5464  (.I0(\edb_top_inst/n2736 ), .I1(\edb_top_inst/n2762 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I3(\edb_top_inst/n2783 ), 
            .O(\edb_top_inst/n2784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5464 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__5465  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .O(\edb_top_inst/n2785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5465 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5466  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/n2785 ), .O(\edb_top_inst/n2786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5466 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5467  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n2787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5467 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5468  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .O(\edb_top_inst/n2788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5468 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5469  (.I0(\edb_top_inst/n2742 ), .I1(\edb_top_inst/n2787 ), 
            .I2(\edb_top_inst/n2788 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .O(\edb_top_inst/n2789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5469 .LUTMASK = 16'h0fee;
    EFX_LUT4 \edb_top_inst/LUT__5470  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I3(\edb_top_inst/la0/la_trig_pos [1]), .O(\edb_top_inst/n2790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5470 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5471  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I1(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n2791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5471 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5472  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [2]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/la0/la_trig_pos [3]), .O(\edb_top_inst/n2792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5472 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5473  (.I0(\edb_top_inst/n2791 ), .I1(\edb_top_inst/la0/la_trig_pos [5]), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), .I3(\edb_top_inst/n2792 ), 
            .O(\edb_top_inst/n2793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5473 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__5474  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .I1(\edb_top_inst/la0/la_trig_pos [8]), .O(\edb_top_inst/n2794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5474 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__5475  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I1(\edb_top_inst/la0/la_trig_pos [4]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I3(\edb_top_inst/la0/la_trig_pos [7]), .O(\edb_top_inst/n2795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5475 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5476  (.I0(\edb_top_inst/n2794 ), .I1(\edb_top_inst/la0/la_trig_pos [6]), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), .I3(\edb_top_inst/n2795 ), 
            .O(\edb_top_inst/n2796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5476 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__5477  (.I0(\edb_top_inst/n2738 ), .I1(\edb_top_inst/n2790 ), 
            .I2(\edb_top_inst/n2793 ), .I3(\edb_top_inst/n2796 ), .O(\edb_top_inst/n2797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5477 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5478  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I2(\edb_top_inst/n2797 ), 
            .I3(\edb_top_inst/n2789 ), .O(\edb_top_inst/n2798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h31ac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5478 .LUTMASK = 16'h31ac;
    EFX_LUT4 \edb_top_inst/LUT__5479  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/n2798 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/n2799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h330e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5479 .LUTMASK = 16'h330e;
    EFX_LUT4 \edb_top_inst/LUT__5480  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/n2763 ), .O(\edb_top_inst/n2800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5480 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5481  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .O(\edb_top_inst/n2801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5481 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5482  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/n2700 ), .I2(\edb_top_inst/n2801 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n2802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5482 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__5483  (.I0(\edb_top_inst/n2784 ), .I1(\edb_top_inst/n2786 ), 
            .I2(\edb_top_inst/n2799 ), .I3(\edb_top_inst/n2802 ), .O(\edb_top_inst/la0/la_biu_inst/next_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5483 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__5484  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), .O(\edb_top_inst/la0/la_biu_inst/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5484 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5485  (.I0(\edb_top_inst/n2079 ), .I1(\edb_top_inst/n2087 ), 
            .I2(\edb_top_inst/n2141 ), .O(\edb_top_inst/n2803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5485 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__5486  (.I0(\edb_top_inst/n2803 ), .I1(\edb_top_inst/n2143 ), 
            .I2(\edb_top_inst/n2144 ), .I3(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5486 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__5487  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), .O(\edb_top_inst/la0/la_biu_inst/n1318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5487 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5488  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5488 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__5489  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/n1902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5489 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5490  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/n2761 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n2804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5490 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__5491  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/n2804 ), 
            .I3(\edb_top_inst/n2763 ), .O(\edb_top_inst/n2805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h73c0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5491 .LUTMASK = 16'h73c0;
    EFX_LUT4 \edb_top_inst/LUT__5492  (.I0(\edb_top_inst/n2773 ), .I1(\edb_top_inst/n2781 ), 
            .O(\edb_top_inst/n2806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5492 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5493  (.I0(\edb_top_inst/n2736 ), .I1(\edb_top_inst/n2762 ), 
            .I2(\edb_top_inst/n2806 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .O(\edb_top_inst/n2807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5493 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__5494  (.I0(\edb_top_inst/n2807 ), .I1(\edb_top_inst/n2785 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I3(\edb_top_inst/n2805 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5494 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__5495  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n19936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5495 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5496  (.I0(\edb_top_inst/n2762 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/n2786 ), .O(\edb_top_inst/n2808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5496 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5497  (.I0(\edb_top_inst/n2781 ), .I1(\edb_top_inst/n2773 ), 
            .I2(\edb_top_inst/n2761 ), .O(\edb_top_inst/n2809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5497 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__5498  (.I0(\edb_top_inst/n2222 ), .I1(\edb_top_inst/n2785 ), 
            .O(\edb_top_inst/n2810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5498 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5499  (.I0(\edb_top_inst/n2809 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/n2763 ), .I3(\edb_top_inst/n2810 ), .O(\edb_top_inst/n2811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5499 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__5500  (.I0(\edb_top_inst/n2801 ), .I1(\edb_top_inst/n2761 ), 
            .I2(\edb_top_inst/n2700 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .O(\edb_top_inst/n2812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5500 .LUTMASK = 16'h77f0;
    EFX_LUT4 \edb_top_inst/LUT__5501  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n2813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5501 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__5502  (.I0(\edb_top_inst/n2812 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .I3(\edb_top_inst/n2813 ), 
            .O(\edb_top_inst/n2814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5502 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__5503  (.I0(\edb_top_inst/n2808 ), .I1(\edb_top_inst/n2736 ), 
            .I2(\edb_top_inst/n2811 ), .I3(\edb_top_inst/n2814 ), .O(\edb_top_inst/la0/la_biu_inst/next_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5503 .LUTMASK = 16'hf2ff;
    EFX_LUT4 \edb_top_inst/LUT__5504  (.I0(\edb_top_inst/n2797 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I3(\edb_top_inst/n2788 ), 
            .O(\edb_top_inst/n2815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5504 .LUTMASK = 16'hec0c;
    EFX_LUT4 \edb_top_inst/LUT__5505  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I2(\edb_top_inst/n2800 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n2816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0dcc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5505 .LUTMASK = 16'h0dcc;
    EFX_LUT4 \edb_top_inst/LUT__5506  (.I0(\edb_top_inst/n2815 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .I3(\edb_top_inst/n2816 ), 
            .O(\edb_top_inst/n2817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7457, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5506 .LUTMASK = 16'h7457;
    EFX_LUT4 \edb_top_inst/LUT__5507  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n2818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5507 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5508  (.I0(\edb_top_inst/n2761 ), .I1(\edb_top_inst/n2742 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .O(\edb_top_inst/n2819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5508 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__5509  (.I0(\edb_top_inst/n2787 ), .I1(\edb_top_inst/n2742 ), 
            .I2(\edb_top_inst/n2797 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .O(\edb_top_inst/n2820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5509 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__5510  (.I0(\edb_top_inst/n2736 ), .I1(\edb_top_inst/n2819 ), 
            .I2(\edb_top_inst/n2820 ), .I3(\edb_top_inst/n2816 ), .O(\edb_top_inst/n2821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5510 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__5511  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/n2806 ), 
            .I2(\edb_top_inst/n2761 ), .I3(\edb_top_inst/n2782 ), .O(\edb_top_inst/n2822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5511 .LUTMASK = 16'hbe00;
    EFX_LUT4 \edb_top_inst/LUT__5512  (.I0(\edb_top_inst/n2822 ), .I1(\edb_top_inst/n2818 ), 
            .I2(\edb_top_inst/n2821 ), .I3(\edb_top_inst/n2817 ), .O(\edb_top_inst/la0/la_biu_inst/next_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c73, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5512 .LUTMASK = 16'h0c73;
    EFX_LUT4 \edb_top_inst/LUT__5513  (.I0(\edb_top_inst/la0/la_biu_inst/n370 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
            .O(\edb_top_inst/ceg_net18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5513 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5514  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5514 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5515  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .O(\edb_top_inst/ceg_net24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5515 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5516  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/n2810 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5516 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__5517  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5517 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__5518  (.I0(\edb_top_inst/la0/la_biu_inst/n1909 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n2823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5518 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5519  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/n2823 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5519 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5520  (.I0(\edb_top_inst/n2788 ), .I1(\edb_top_inst/n2222 ), 
            .I2(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5520 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__5521  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5521 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5522  (.I0(\edb_top_inst/n2823 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/~ceg_net27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5522 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5523  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n2223 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5523 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__5524  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [15]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5524 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5525  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [16]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5525 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5526  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [17]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5526 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5527  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [18]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5527 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5528  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [19]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5528 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5529  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [5]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [20]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5529 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5530  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [21]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5530 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5531  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [7]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [22]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5531 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5532  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [23]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5532 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5533  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [24]), .I2(\edb_top_inst/n2223 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5533 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5534  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), 
            .I1(\edb_top_inst/n2681 ), .O(\edb_top_inst/n2824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5534 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5535  (.I0(\edb_top_inst/n2693 ), .I1(\edb_top_inst/n2824 ), 
            .O(\edb_top_inst/n2825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5535 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5536  (.I0(\edb_top_inst/n2717 ), .I1(\edb_top_inst/n2732 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
            .I3(\edb_top_inst/n2825 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5536 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__5537  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/n2683 ), .O(\edb_top_inst/n2826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5537 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5538  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .I2(\edb_top_inst/la0/la_window_depth [0]), 
            .O(\edb_top_inst/n2827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5538 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5539  (.I0(\edb_top_inst/n2827 ), .I1(\edb_top_inst/n2707 ), 
            .O(\edb_top_inst/n2828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5539 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5540  (.I0(\edb_top_inst/n2826 ), .I1(\edb_top_inst/n2687 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1]), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5540 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5541  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n2685 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n2829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h010e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5541 .LUTMASK = 16'h010e;
    EFX_LUT4 \edb_top_inst/LUT__5542  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5542 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5543  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), .I2(\edb_top_inst/n2830 ), 
            .I3(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5543 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__5544  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n2693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2]), 
            .I3(\edb_top_inst/n2829 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5544 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5545  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/la0/la_window_depth [4]), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0130, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5545 .LUTMASK = 16'h0130;
    EFX_LUT4 \edb_top_inst/LUT__5546  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), .I2(\edb_top_inst/la0/la_window_depth [0]), 
            .O(\edb_top_inst/n2833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5546 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5547  (.I0(\edb_top_inst/n2833 ), .I1(\edb_top_inst/n2827 ), 
            .I2(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n2834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5547 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5548  (.I0(\edb_top_inst/n2834 ), .I1(\edb_top_inst/n2693 ), 
            .O(\edb_top_inst/n2835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5548 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5549  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3]), 
            .I1(\edb_top_inst/n2832 ), .I2(\edb_top_inst/n2835 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5549 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5550  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .O(\edb_top_inst/n2836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5550 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5551  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/n2836 ), .O(\edb_top_inst/n2837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5551 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5552  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5552 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5553  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5553 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5554  (.I0(\edb_top_inst/n2839 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5554 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5555  (.I0(\edb_top_inst/n2840 ), .I1(\edb_top_inst/n2824 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n2679 ), 
            .O(\edb_top_inst/n2841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5555 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__5556  (.I0(\edb_top_inst/n2837 ), .I1(\edb_top_inst/n2832 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4]), 
            .I3(\edb_top_inst/n2841 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5556 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5557  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/n2827 ), .O(\edb_top_inst/n2842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5557 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5558  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5558 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5559  (.I0(\edb_top_inst/n2843 ), .I1(\edb_top_inst/n2839 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5559 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5560  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/n2842 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n2679 ), 
            .O(\edb_top_inst/n2845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5560 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__5561  (.I0(\edb_top_inst/n2836 ), .I1(\edb_top_inst/n2832 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5]), 
            .I3(\edb_top_inst/n2845 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5561 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5562  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/n2685 ), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n2846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5562 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__5563  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5563 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5564  (.I0(\edb_top_inst/n2847 ), .I1(\edb_top_inst/n2843 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5564 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5565  (.I0(\edb_top_inst/n2848 ), .I1(\edb_top_inst/n2831 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n2679 ), 
            .O(\edb_top_inst/n2849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5565 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__5566  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6]), 
            .I1(\edb_top_inst/n2846 ), .I2(\edb_top_inst/n2849 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5566 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5567  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5567 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5568  (.I0(\edb_top_inst/n2850 ), .I1(\edb_top_inst/n2847 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5568 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5569  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2834 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n2679 ), 
            .O(\edb_top_inst/n2852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5569 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__5570  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/n2718 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7]), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5570 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5571  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/n2718 ), 
            .O(\edb_top_inst/n2853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5571 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__5572  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5572 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5573  (.I0(\edb_top_inst/n2854 ), .I1(\edb_top_inst/n2850 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5573 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5574  (.I0(\edb_top_inst/n2855 ), .I1(\edb_top_inst/n2824 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5574 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__5575  (.I0(\edb_top_inst/n2840 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/n2856 ), 
            .O(\edb_top_inst/n2857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5575 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__5576  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8]), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5576 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5577  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5577 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5578  (.I0(\edb_top_inst/n2858 ), .I1(\edb_top_inst/n2854 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5578 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5579  (.I0(\edb_top_inst/n2859 ), .I1(\edb_top_inst/n2842 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5579 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__5580  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/n2860 ), 
            .O(\edb_top_inst/n2861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5580 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__5581  (.I0(\edb_top_inst/n2732 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9]), 
            .I2(\edb_top_inst/n2861 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5581 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5582  (.I0(\edb_top_inst/n2717 ), .I1(\edb_top_inst/n2732 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
            .I3(\edb_top_inst/n2825 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5582 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__5583  (.I0(\edb_top_inst/n2826 ), .I1(\edb_top_inst/n2687 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1]), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5583 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5584  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n2693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2]), 
            .I3(\edb_top_inst/n2829 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5584 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5585  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3]), 
            .I1(\edb_top_inst/n2832 ), .I2(\edb_top_inst/n2835 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5585 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5586  (.I0(\edb_top_inst/n2837 ), .I1(\edb_top_inst/n2832 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4]), 
            .I3(\edb_top_inst/n2841 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5586 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5587  (.I0(\edb_top_inst/n2836 ), .I1(\edb_top_inst/n2832 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5]), 
            .I3(\edb_top_inst/n2845 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5587 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5588  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6]), 
            .I1(\edb_top_inst/n2846 ), .I2(\edb_top_inst/n2849 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5588 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5589  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/n2718 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7]), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5589 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5590  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8]), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5590 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5591  (.I0(\edb_top_inst/n2732 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9]), 
            .I2(\edb_top_inst/n2861 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5591 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5592  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [3]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [1]), .O(\edb_top_inst/la0/n617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5592 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5593  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/la0/module_state [2]), 
            .I3(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n2862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5593 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__5594  (.I0(\edb_top_inst/n2862 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr [81]), .I3(jtag_inst1_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5594 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5595  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5595 .LUTMASK = 16'h8888;
    EFX_ADD \edb_top_inst/la0/add_1054/i1  (.I0(\edb_top_inst/la0/address_counter [16]), 
            .I1(\edb_top_inst/la0/address_counter [15]), .CI(1'b0), .O(\edb_top_inst/la0/n1818 [1]), 
            .CO(\edb_top_inst/la0/add_1054/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i1  (.I0(\edb_top_inst/la0/address_counter [0]), 
            .I1(\edb_top_inst/la0/n616 ), .CI(1'b0), .O(\edb_top_inst/la0/n1837 [0]), 
            .CO(\edb_top_inst/la0/add_98/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1057/i1  (.I0(\edb_top_inst/la0/bit_count [1]), 
            .I1(\edb_top_inst/la0/bit_count [0]), .CI(1'b0), .O(\edb_top_inst/la0/n1984 [1]), 
            .CO(\edb_top_inst/la0/add_1057/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/add_1057/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1057/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i1  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/trigger_skipper_n/n73 [1]), 
            .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(1'b1), .CI(n2835), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10  (.I0(\edb_top_inst/la0/la_sample_cnt [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9  (.I0(\edb_top_inst/la0/la_sample_cnt [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [9]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8  (.I0(\edb_top_inst/la0/la_sample_cnt [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7  (.I0(\edb_top_inst/la0/la_sample_cnt [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6  (.I0(\edb_top_inst/la0/la_sample_cnt [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5  (.I0(\edb_top_inst/la0/la_sample_cnt [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4  (.I0(\edb_top_inst/la0/la_sample_cnt [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3  (.I0(\edb_top_inst/la0/la_sample_cnt [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [9]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4685)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i63  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n124 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i63 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i63 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i62  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n122 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [62]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i62 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i62 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i61  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n120 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [61]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i61 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i61 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i60  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n118 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [60]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i60 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i60 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), .CI(1'b0), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4696)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(\edb_top_inst/la0/la_sample_cnt [0]), .CI(1'b0), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4710)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .CI(1'b0), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i59  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n116 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [59]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i59 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i59 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i58  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n114 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [58]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i58 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i58 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i57  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n112 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [57]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i57 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i57 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i56  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n110 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [56]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i56 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i56 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i55  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n108 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [55]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i55 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i55 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i54  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n106 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [54]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i54 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i54 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i53  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n104 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [53]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i53 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i53 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i52  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n102 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [52]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i52 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i52 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i51  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n100 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [51]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i51 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i51 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i50  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n98 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [50]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i50 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i50 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i49  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n96 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [49]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i49 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i49 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i48  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n94 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [48]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i48 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i48 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i47  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n92 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [47]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i47 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i47 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i46  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n90 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [46]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i46 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i46 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i45  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n88 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [45]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i45 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i45 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i44  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n86 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [44]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i44 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i44 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i43  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n84 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [43]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i43 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i43 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i42  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n82 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [42]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i42 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i42 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i41  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n80 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [41]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i41 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i41 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i40  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n78 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [40]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i40 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i40 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i39  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n76 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [39]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i39 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i39 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i38  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n74 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [38]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i38 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i38 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i37  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n72 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [37]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i37 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i37 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i36  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n70 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [36]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i36 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i36 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i35  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n68 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [35]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i35 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i35 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i34  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n66 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [34]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i34 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i34 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i33  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n64 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [33]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i33 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i33 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i32  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n62 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [32]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i32 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i31  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n60 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [31]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i31 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i30  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n58 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [30]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i30 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i29  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n56 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [29]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i29 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i28  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n54 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [28]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i28 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i27  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n52 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [27]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i26  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n50 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [26]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i25  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n48 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [25]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i24  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n46 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [24]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i23  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n44 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [23]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i22  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n42 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [22]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i21  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n40 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [21]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i20  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n38 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [20]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i19  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n36 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [19]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i18  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n34 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [18]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i17  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n32 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [17]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i16  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n30 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [16]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i15  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n28 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [15]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i14  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n26 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [14]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i13  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n24 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [13]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i12  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n22 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [12]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i11  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n20 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [11]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i10  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n18 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [10]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i9  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n16 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [9]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i8  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n14 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [8]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i7  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n12 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [7]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i6  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n10 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [6]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i5  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n8 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [5]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i4  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n6 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [4]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i3  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n4 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [3]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i2  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n2 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [2]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5878)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1057/i5  (.I0(\edb_top_inst/la0/bit_count [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1057/n8 ), .O(\edb_top_inst/la0/n1984 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/add_1057/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1057/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1057/i4  (.I0(\edb_top_inst/la0/bit_count [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1057/n6 ), .O(\edb_top_inst/la0/n1984 [4]), 
            .CO(\edb_top_inst/la0/add_1057/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/add_1057/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1057/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1057/i3  (.I0(\edb_top_inst/la0/bit_count [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1057/n4 ), .O(\edb_top_inst/la0/n1984 [3]), 
            .CO(\edb_top_inst/la0/add_1057/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/add_1057/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1057/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1057/i2  (.I0(\edb_top_inst/la0/bit_count [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1057/n2 ), .O(\edb_top_inst/la0/n1984 [2]), 
            .CO(\edb_top_inst/la0/add_1057/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3745)
    defparam \edb_top_inst/la0/add_1057/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1057/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i25  (.I0(\edb_top_inst/la0/address_counter [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n48 ), .O(\edb_top_inst/la0/n1837 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i24  (.I0(\edb_top_inst/la0/address_counter [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n46 ), .O(\edb_top_inst/la0/n1837 [23]), 
            .CO(\edb_top_inst/la0/add_98/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i23  (.I0(\edb_top_inst/la0/address_counter [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n44 ), .O(\edb_top_inst/la0/n1837 [22]), 
            .CO(\edb_top_inst/la0/add_98/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i22  (.I0(\edb_top_inst/la0/address_counter [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n42 ), .O(\edb_top_inst/la0/n1837 [21]), 
            .CO(\edb_top_inst/la0/add_98/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i21  (.I0(\edb_top_inst/la0/address_counter [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n40 ), .O(\edb_top_inst/la0/n1837 [20]), 
            .CO(\edb_top_inst/la0/add_98/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i20  (.I0(\edb_top_inst/la0/address_counter [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n38 ), .O(\edb_top_inst/la0/n1837 [19]), 
            .CO(\edb_top_inst/la0/add_98/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i19  (.I0(\edb_top_inst/la0/address_counter [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n36 ), .O(\edb_top_inst/la0/n1837 [18]), 
            .CO(\edb_top_inst/la0/add_98/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i18  (.I0(\edb_top_inst/la0/address_counter [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n34 ), .O(\edb_top_inst/la0/n1837 [17]), 
            .CO(\edb_top_inst/la0/add_98/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i17  (.I0(\edb_top_inst/la0/address_counter [16]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n32 ), .O(\edb_top_inst/la0/n1837 [16]), 
            .CO(\edb_top_inst/la0/add_98/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i16  (.I0(\edb_top_inst/la0/address_counter [15]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n30 ), .O(\edb_top_inst/la0/n1837 [15]), 
            .CO(\edb_top_inst/la0/add_98/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i15  (.I0(\edb_top_inst/la0/address_counter [14]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n28 ), .O(\edb_top_inst/la0/n1837 [14]), 
            .CO(\edb_top_inst/la0/add_98/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i14  (.I0(\edb_top_inst/la0/address_counter [13]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n26 ), .O(\edb_top_inst/la0/n1837 [13]), 
            .CO(\edb_top_inst/la0/add_98/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i13  (.I0(\edb_top_inst/la0/address_counter [12]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n24 ), .O(\edb_top_inst/la0/n1837 [12]), 
            .CO(\edb_top_inst/la0/add_98/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i12  (.I0(\edb_top_inst/la0/address_counter [11]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n22 ), .O(\edb_top_inst/la0/n1837 [11]), 
            .CO(\edb_top_inst/la0/add_98/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i11  (.I0(\edb_top_inst/la0/address_counter [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n20 ), .O(\edb_top_inst/la0/n1837 [10]), 
            .CO(\edb_top_inst/la0/add_98/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i10  (.I0(\edb_top_inst/la0/address_counter [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n18 ), .O(\edb_top_inst/la0/n1837 [9]), 
            .CO(\edb_top_inst/la0/add_98/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i9  (.I0(\edb_top_inst/la0/address_counter [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n16 ), .O(\edb_top_inst/la0/n1837 [8]), 
            .CO(\edb_top_inst/la0/add_98/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i8  (.I0(\edb_top_inst/la0/address_counter [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n14 ), .O(\edb_top_inst/la0/n1837 [7]), 
            .CO(\edb_top_inst/la0/add_98/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i7  (.I0(\edb_top_inst/la0/address_counter [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n12 ), .O(\edb_top_inst/la0/n1837 [6]), 
            .CO(\edb_top_inst/la0/add_98/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i6  (.I0(\edb_top_inst/la0/address_counter [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n10 ), .O(\edb_top_inst/la0/n1837 [5]), 
            .CO(\edb_top_inst/la0/add_98/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i5  (.I0(\edb_top_inst/la0/address_counter [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n8 ), .O(\edb_top_inst/la0/n1837 [4]), 
            .CO(\edb_top_inst/la0/add_98/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i4  (.I0(\edb_top_inst/la0/address_counter [3]), 
            .I1(\edb_top_inst/la0/n619 ), .CI(\edb_top_inst/la0/add_98/n6 ), 
            .O(\edb_top_inst/la0/n1837 [3]), .CO(\edb_top_inst/la0/add_98/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i3  (.I0(\edb_top_inst/la0/address_counter [2]), 
            .I1(\edb_top_inst/la0/n618 ), .CI(\edb_top_inst/la0/add_98/n4 ), 
            .O(\edb_top_inst/la0/n1837 [2]), .CO(\edb_top_inst/la0/add_98/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i2  (.I0(\edb_top_inst/la0/address_counter [1]), 
            .I1(\edb_top_inst/la0/n617 ), .CI(\edb_top_inst/la0/add_98/n2 ), 
            .O(\edb_top_inst/la0/n1837 [1]), .CO(\edb_top_inst/la0/add_98/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3718)
    defparam \edb_top_inst/la0/add_98/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i9  (.I0(\edb_top_inst/la0/address_counter [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n16 ), .O(\edb_top_inst/la0/n1818 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i8  (.I0(\edb_top_inst/la0/address_counter [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n14 ), .O(\edb_top_inst/la0/n1818 [8]), 
            .CO(\edb_top_inst/la0/add_1054/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i7  (.I0(\edb_top_inst/la0/address_counter [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n12 ), .O(\edb_top_inst/la0/n1818 [7]), 
            .CO(\edb_top_inst/la0/add_1054/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i6  (.I0(\edb_top_inst/la0/address_counter [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n10 ), .O(\edb_top_inst/la0/n1818 [6]), 
            .CO(\edb_top_inst/la0/add_1054/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i5  (.I0(\edb_top_inst/la0/address_counter [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n8 ), .O(\edb_top_inst/la0/n1818 [5]), 
            .CO(\edb_top_inst/la0/add_1054/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i4  (.I0(\edb_top_inst/la0/address_counter [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n6 ), .O(\edb_top_inst/la0/n1818 [4]), 
            .CO(\edb_top_inst/la0/add_1054/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i3  (.I0(\edb_top_inst/la0/address_counter [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n4 ), .O(\edb_top_inst/la0/n1818 [3]), 
            .CO(\edb_top_inst/la0/add_1054/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1054/i2  (.I0(\edb_top_inst/la0/address_counter [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1054/n2 ), .O(\edb_top_inst/la0/n1818 [2]), 
            .CO(\edb_top_inst/la0/add_1054/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3717)
    defparam \edb_top_inst/la0/add_1054/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1054/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [29:25]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [29:25]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [24:23], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [1], 
            2'b00}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [24:20]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [14], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [37:35]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [39:35]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [14:13], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [0], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [11:10]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [14:10]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [34:30]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [34:30]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [9], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [29:26]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [9:5]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [18], 
            3'b000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [19:15]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [25:23], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [1:0]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [4:0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n646 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [44:43], 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [18], 
            2'b00}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [44:40]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(454)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h1 .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__8044 (.I0(b[0]), .I1(a[0]), .O(n26[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(35)
    defparam LUT__8044.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8045 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [4]), 
            .O(rx_data[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8045.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8046 (.I0(\uart_rx_inst/r_Clock_Count [3]), .I1(\uart_rx_inst/r_Clock_Count [6]), 
            .O(n2768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8046.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8047 (.I0(\uart_rx_inst/r_Clock_Count [1]), .I1(\uart_rx_inst/r_Clock_Count [0]), 
            .I2(\uart_rx_inst/r_Clock_Count [2]), .O(n2769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__8047.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__8048 (.I0(\uart_rx_inst/r_Clock_Count [5]), .I1(\uart_rx_inst/r_Clock_Count [4]), 
            .I2(\uart_rx_inst/r_Clock_Count [6]), .O(n2770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__8048.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__8049 (.I0(\uart_rx_inst/r_Clock_Count [7]), .I1(\uart_rx_inst/r_Clock_Count [8]), 
            .O(n2771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8049.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8050 (.I0(n2769), .I1(n2768), .I2(n2770), .I3(n2771), 
            .O(n2772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__8050.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__8051 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(\uart_rx_inst/r_Clock_Count [16]), 
            .I2(\uart_rx_inst/r_Clock_Count [20]), .I3(\uart_rx_inst/r_Clock_Count [22]), 
            .O(n2773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8051.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8052 (.I0(\uart_rx_inst/r_Clock_Count [13]), .I1(\uart_rx_inst/r_Clock_Count [15]), 
            .I2(\uart_rx_inst/r_Clock_Count [19]), .O(n2774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8052.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8053 (.I0(n2773), .I1(n2774), .O(n2775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8053.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8054 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(\uart_rx_inst/r_Clock_Count [29]), 
            .I2(\uart_rx_inst/r_Clock_Count [30]), .I3(\uart_rx_inst/r_Clock_Count [31]), 
            .O(n2776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8054.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8055 (.I0(\uart_rx_inst/r_Clock_Count [24]), .I1(\uart_rx_inst/r_Clock_Count [25]), 
            .I2(\uart_rx_inst/r_Clock_Count [26]), .I3(\uart_rx_inst/r_Clock_Count [27]), 
            .O(n2777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8055.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8056 (.I0(\uart_rx_inst/r_Clock_Count [17]), .I1(\uart_rx_inst/r_Clock_Count [18]), 
            .I2(\uart_rx_inst/r_Clock_Count [21]), .I3(\uart_rx_inst/r_Clock_Count [23]), 
            .O(n2778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8056.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8057 (.I0(\uart_rx_inst/r_Clock_Count [9]), .I1(\uart_rx_inst/r_Clock_Count [10]), 
            .I2(\uart_rx_inst/r_Clock_Count [11]), .I3(\uart_rx_inst/r_Clock_Count [12]), 
            .O(n2779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8057.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8058 (.I0(n2776), .I1(n2777), .I2(n2778), .I3(n2779), 
            .O(n2780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8058.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8059 (.I0(\uart_rx_inst/r_SM_Main [2]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .O(\uart_rx_inst/n924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8059.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8060 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/n924 ), 
            .O(n2781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8060.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8061 (.I0(n2772), .I1(n2780), .I2(n2775), .I3(n2781), 
            .O(n2782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__8061.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__8062 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(n2782), .O(\uart_rx_inst/n925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8062.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8063 (.I0(n2772), .I1(n2775), .I2(n2780), .O(\uart_rx_inst/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(137)
    defparam LUT__8063.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__8064 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .O(n2783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8064.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8065 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(n2783), .O(n2784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__8065.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8066 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [2]), 
            .I2(\uart_rx_inst/r_Clock_Count [3]), .I3(\uart_rx_inst/r_Clock_Count [4]), 
            .O(n2785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__8066.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8067 (.I0(\uart_rx_inst/r_Clock_Count [5]), .I1(\uart_rx_inst/r_Clock_Count [8]), 
            .I2(\uart_rx_inst/r_Clock_Count [1]), .O(n2786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8067.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8068 (.I0(\uart_rx_inst/r_Clock_Count [6]), .I1(\uart_rx_inst/r_Clock_Count [7]), 
            .I2(n2785), .I3(n2786), .O(n2787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8068.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8069 (.I0(\uart_rx_inst/r_SM_Main [1]), .I1(\uart_rx_inst/r_SM_Main [0]), 
            .O(n2788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8069.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8070 (.I0(n2787), .I1(n2780), .I2(n2775), .I3(n2788), 
            .O(n2789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__8070.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__8071 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(n2773), .I3(n2774), .O(n2790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8071.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8072 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(\uart_rx_inst/r_Rx_Data ), .O(n2791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8072.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8073 (.I0(n2772), .I1(n2780), .I2(n2790), .I3(n2791), 
            .O(n2792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__8073.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__8074 (.I0(n2784), .I1(\uart_rx_inst/n151 ), .I2(n2789), 
            .I3(n2792), .O(\uart_rx_inst/n896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8074.LUTMASK = 16'hf2ff;
    EFX_LUT4 LUT__8075 (.I0(n2772), .I1(\uart_rx_inst/r_SM_Main [1]), .I2(n2775), 
            .I3(n2780), .O(n2793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__8075.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8076 (.I0(n2793), .I1(n2789), .I2(\uart_rx_inst/r_Clock_Count [0]), 
            .O(\uart_rx_inst/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8076.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__8077 (.I0(\uart_rx_inst/r_Rx_Data ), .I1(n2789), .I2(n2788), 
            .I3(\uart_rx_inst/r_SM_Main [2]), .O(ceg_net14)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(88)
    defparam LUT__8077.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__8078 (.I0(\uart_rx_inst/r_SM_Main [2]), .I1(\uart_rx_inst/n151 ), 
            .I2(\uart_rx_inst/r_SM_Main [0]), .I3(\uart_rx_inst/r_SM_Main [1]), 
            .O(ceg_net32)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(88)
    defparam LUT__8078.LUTMASK = 16'heff0;
    EFX_LUT4 LUT__8079 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .O(\uart_rx_inst/n903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(151)
    defparam LUT__8079.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8080 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_SM_Main [2]), 
            .I2(n2793), .O(ceg_net26)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(88)
    defparam LUT__8080.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__8081 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(\uart_rx_inst/r_Bit_Index [0]), .I3(n2782), .O(\uart_rx_inst/n959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8081.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8082 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(\uart_rx_inst/r_Bit_Index [1]), .I3(n2782), .O(\uart_rx_inst/n961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8082.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8083 (.I0(\uart_rx_inst/r_Bit_Index [2]), .I1(n2782), 
            .I2(n2783), .O(\uart_rx_inst/n963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8083.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__8084 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(n2782), .O(\uart_rx_inst/n965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8084.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8085 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(\uart_rx_inst/r_Bit_Index [0]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(n2782), .O(\uart_rx_inst/n967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8085.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8086 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(n2782), .O(\uart_rx_inst/n969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8086.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8087 (.I0(\uart_rx_inst/r_Bit_Index [2]), .I1(n2782), 
            .I2(n2783), .O(\uart_rx_inst/n971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8087.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8088 (.I0(\uart_rx_inst/r_Rx_Data ), .I1(n2780), .I2(n2775), 
            .I3(n2787), .O(n2794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8088.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8089 (.I0(n2794), .I1(\uart_rx_inst/n151 ), .I2(\uart_rx_inst/r_SM_Main [0]), 
            .I3(\uart_rx_inst/r_SM_Main [1]), .O(\uart_rx_inst/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfa0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8089.LUTMASK = 16'hcfa0;
    EFX_LUT4 LUT__8090 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/n924 ), 
            .O(\uart_rx_inst/n955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(17)
    defparam LUT__8090.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8091 (.I0(n2789), .I1(n2793), .I2(\uart_rx_inst/r_Clock_Count [0]), 
            .I3(\uart_rx_inst/r_Clock_Count [1]), .O(\uart_rx_inst/n767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8091.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__8092 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [1]), 
            .O(n2795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8092.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8093 (.I0(n2789), .I1(n2793), .I2(\uart_rx_inst/r_Clock_Count [2]), 
            .I3(n2795), .O(\uart_rx_inst/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8093.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__8094 (.I0(\uart_rx_inst/r_Clock_Count [2]), .I1(n2795), 
            .I2(\uart_rx_inst/r_Clock_Count [3]), .O(n2796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__8094.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__8095 (.I0(n2793), .I1(n2789), .I2(n2796), .O(\uart_rx_inst/n773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8095.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__8096 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [1]), 
            .I2(\uart_rx_inst/r_Clock_Count [2]), .I3(\uart_rx_inst/r_Clock_Count [3]), 
            .O(n2797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8096.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8097 (.I0(n2789), .I1(n2793), .I2(\uart_rx_inst/r_Clock_Count [4]), 
            .I3(n2797), .O(\uart_rx_inst/n776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8097.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__8098 (.I0(\uart_rx_inst/r_Clock_Count [4]), .I1(n2797), 
            .O(n2798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8098.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8099 (.I0(n2789), .I1(n2793), .I2(\uart_rx_inst/r_Clock_Count [5]), 
            .I3(n2798), .O(\uart_rx_inst/n779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8099.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__8100 (.I0(\uart_rx_inst/r_Clock_Count [5]), .I1(n2798), 
            .I2(\uart_rx_inst/r_Clock_Count [6]), .O(n2799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__8100.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__8101 (.I0(n2793), .I1(n2789), .I2(n2799), .O(\uart_rx_inst/n782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8101.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__8102 (.I0(\uart_rx_inst/r_Clock_Count [5]), .I1(\uart_rx_inst/r_Clock_Count [6]), 
            .I2(n2798), .I3(\uart_rx_inst/r_Clock_Count [7]), .O(n2800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__8102.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__8103 (.I0(n2793), .I1(n2789), .I2(n2800), .O(\uart_rx_inst/n785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8103.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__8104 (.I0(\uart_rx_inst/r_Clock_Count [4]), .I1(\uart_rx_inst/r_Clock_Count [5]), 
            .I2(\uart_rx_inst/r_Clock_Count [6]), .I3(\uart_rx_inst/r_Clock_Count [7]), 
            .O(n2801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8104.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8105 (.I0(n2797), .I1(n2801), .O(n2802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8105.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8106 (.I0(n2789), .I1(n2793), .I2(\uart_rx_inst/r_Clock_Count [8]), 
            .I3(n2802), .O(\uart_rx_inst/n788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8106.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__8107 (.I0(\uart_rx_inst/r_Clock_Count [8]), .I1(n2802), 
            .I2(\uart_rx_inst/r_Clock_Count [9]), .I3(n2789), .O(\uart_rx_inst/n791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8107.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8108 (.I0(\uart_rx_inst/r_Clock_Count [8]), .I1(\uart_rx_inst/r_Clock_Count [9]), 
            .I2(n2802), .O(n2803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8108.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8109 (.I0(\uart_rx_inst/r_Clock_Count [10]), .I1(n2803), 
            .I2(n2789), .O(\uart_rx_inst/n794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8109.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8110 (.I0(\uart_rx_inst/r_Clock_Count [10]), .I1(n2803), 
            .I2(\uart_rx_inst/r_Clock_Count [11]), .I3(n2789), .O(\uart_rx_inst/n797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8110.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8111 (.I0(\uart_rx_inst/r_Clock_Count [8]), .I1(\uart_rx_inst/r_Clock_Count [9]), 
            .I2(\uart_rx_inst/r_Clock_Count [10]), .I3(\uart_rx_inst/r_Clock_Count [11]), 
            .O(n2804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8111.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8112 (.I0(n2797), .I1(n2801), .I2(n2804), .O(n2805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8112.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8113 (.I0(\uart_rx_inst/r_Clock_Count [12]), .I1(n2805), 
            .I2(n2789), .O(\uart_rx_inst/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8113.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8114 (.I0(\uart_rx_inst/r_Clock_Count [12]), .I1(n2805), 
            .I2(\uart_rx_inst/r_Clock_Count [13]), .I3(n2789), .O(\uart_rx_inst/n803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8114.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8115 (.I0(\uart_rx_inst/r_Clock_Count [12]), .I1(\uart_rx_inst/r_Clock_Count [13]), 
            .O(n2806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8115.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8116 (.I0(n2797), .I1(n2801), .I2(n2804), .I3(n2806), 
            .O(n2807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8116.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8117 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(n2807), 
            .I2(n2789), .O(\uart_rx_inst/n806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8117.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8118 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(n2807), 
            .O(n2808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8118.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8119 (.I0(\uart_rx_inst/r_Clock_Count [15]), .I1(n2808), 
            .I2(n2789), .O(\uart_rx_inst/n809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8119.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8120 (.I0(\uart_rx_inst/r_Clock_Count [15]), .I1(n2808), 
            .I2(\uart_rx_inst/r_Clock_Count [16]), .I3(n2789), .O(\uart_rx_inst/n812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8120.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8121 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(\uart_rx_inst/r_Clock_Count [15]), 
            .I2(\uart_rx_inst/r_Clock_Count [16]), .O(n2809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8121.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8122 (.I0(n2807), .I1(n2809), .I2(\uart_rx_inst/r_Clock_Count [17]), 
            .I3(n2789), .O(\uart_rx_inst/n815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8122.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8123 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(\uart_rx_inst/r_Clock_Count [15]), 
            .I2(\uart_rx_inst/r_Clock_Count [16]), .I3(\uart_rx_inst/r_Clock_Count [17]), 
            .O(n2810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8123.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8124 (.I0(n2805), .I1(n2806), .I2(n2810), .O(n2811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8124.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8125 (.I0(\uart_rx_inst/r_Clock_Count [18]), .I1(n2811), 
            .I2(n2789), .O(\uart_rx_inst/n818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8125.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8126 (.I0(\uart_rx_inst/r_Clock_Count [18]), .I1(n2811), 
            .I2(\uart_rx_inst/r_Clock_Count [19]), .I3(n2789), .O(\uart_rx_inst/n821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8126.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8127 (.I0(\uart_rx_inst/r_Clock_Count [18]), .I1(\uart_rx_inst/r_Clock_Count [19]), 
            .O(n2812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8127.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8128 (.I0(n2807), .I1(n2810), .I2(n2812), .O(n2813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8128.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8129 (.I0(\uart_rx_inst/r_Clock_Count [20]), .I1(n2813), 
            .I2(n2789), .O(\uart_rx_inst/n824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8129.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8130 (.I0(\uart_rx_inst/r_Clock_Count [20]), .I1(n2813), 
            .I2(\uart_rx_inst/r_Clock_Count [21]), .I3(n2789), .O(\uart_rx_inst/n827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8130.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8131 (.I0(\uart_rx_inst/r_Clock_Count [18]), .I1(\uart_rx_inst/r_Clock_Count [19]), 
            .I2(\uart_rx_inst/r_Clock_Count [20]), .I3(\uart_rx_inst/r_Clock_Count [21]), 
            .O(n2814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8131.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8132 (.I0(n2807), .I1(n2810), .I2(n2814), .O(n2815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8132.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8133 (.I0(\uart_rx_inst/r_Clock_Count [22]), .I1(n2815), 
            .I2(n2789), .O(\uart_rx_inst/n830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8133.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8134 (.I0(\uart_rx_inst/r_Clock_Count [22]), .I1(n2815), 
            .I2(\uart_rx_inst/r_Clock_Count [23]), .I3(n2789), .O(\uart_rx_inst/n833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8134.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8135 (.I0(\uart_rx_inst/r_Clock_Count [22]), .I1(\uart_rx_inst/r_Clock_Count [23]), 
            .O(n2816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8135.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8136 (.I0(n2815), .I1(n2816), .I2(\uart_rx_inst/r_Clock_Count [24]), 
            .I3(n2789), .O(\uart_rx_inst/n836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8136.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8137 (.I0(\uart_rx_inst/r_Clock_Count [22]), .I1(\uart_rx_inst/r_Clock_Count [23]), 
            .I2(\uart_rx_inst/r_Clock_Count [24]), .O(n2817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8137.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8138 (.I0(n2815), .I1(n2817), .I2(\uart_rx_inst/r_Clock_Count [25]), 
            .I3(n2789), .O(\uart_rx_inst/n839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8138.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8139 (.I0(\uart_rx_inst/r_Clock_Count [25]), .I1(n2810), 
            .I2(n2814), .I3(n2817), .O(n2818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8139.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8140 (.I0(n2807), .I1(n2818), .O(n2819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8140.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8141 (.I0(\uart_rx_inst/r_Clock_Count [26]), .I1(n2819), 
            .I2(n2789), .O(\uart_rx_inst/n842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8141.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8142 (.I0(\uart_rx_inst/r_Clock_Count [26]), .I1(n2819), 
            .I2(\uart_rx_inst/r_Clock_Count [27]), .I3(n2789), .O(\uart_rx_inst/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8142.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8143 (.I0(\uart_rx_inst/r_Clock_Count [26]), .I1(\uart_rx_inst/r_Clock_Count [27]), 
            .I2(n2807), .I3(n2818), .O(n2820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8143.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8144 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(n2820), 
            .I2(n2789), .O(\uart_rx_inst/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8144.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8145 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(n2820), 
            .I2(\uart_rx_inst/r_Clock_Count [29]), .I3(n2789), .O(\uart_rx_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8145.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8146 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(\uart_rx_inst/r_Clock_Count [29]), 
            .O(n2821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8146.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8147 (.I0(n2820), .I1(n2821), .I2(\uart_rx_inst/r_Clock_Count [30]), 
            .I3(n2789), .O(\uart_rx_inst/n854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8147.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8148 (.I0(\uart_rx_inst/r_Clock_Count [30]), .I1(n2821), 
            .O(n2822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8148.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8149 (.I0(n2820), .I1(n2822), .I2(\uart_rx_inst/r_Clock_Count [31]), 
            .I3(n2789), .O(\uart_rx_inst/n857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(175)
    defparam LUT__8149.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8150 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_SM_Main [1]), .O(\uart_rx_inst/n861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(151)
    defparam LUT__8150.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8151 (.I0(\uart_rx_inst/r_Bit_Index [2]), .I1(n2783), 
            .I2(\uart_rx_inst/r_SM_Main [1]), .O(\uart_rx_inst/n865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(151)
    defparam LUT__8151.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8152 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [1]), 
            .O(rx_data[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8152.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8153 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [2]), 
            .O(rx_data[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8153.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8154 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [3]), 
            .O(rx_data[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8154.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8155 (.I0(\uart_tx_inst/r_Clock_Count [1]), .I1(\uart_tx_inst/r_Clock_Count [0]), 
            .I2(\uart_tx_inst/r_Clock_Count [2]), .I3(\uart_tx_inst/r_Clock_Count [3]), 
            .O(n2823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__8155.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__8156 (.I0(\uart_tx_inst/r_Clock_Count [4]), .I1(\uart_tx_inst/r_Clock_Count [5]), 
            .O(n2824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8156.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8157 (.I0(\uart_tx_inst/r_Clock_Count [7]), .I1(\uart_tx_inst/r_Clock_Count [8]), 
            .O(n2825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8157.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8158 (.I0(n2823), .I1(n2824), .I2(\uart_tx_inst/r_Clock_Count [6]), 
            .I3(n2825), .O(\uart_tx_inst/LessThan_9/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bff */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(242)
    defparam LUT__8158.LUTMASK = 16'h0bff;
    EFX_LUT4 LUT__8159 (.I0(\uart_tx_inst/r_SM_Main [1]), .I1(\uart_tx_inst/r_SM_Main [0]), 
            .I2(\uart_tx_inst/LessThan_9/n18 ), .O(n2826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__8159.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__8160 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(n2826), 
            .O(\uart_tx_inst/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8160.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8161 (.I0(\uart_tx_inst/r_Tx_Data [4]), .I1(\uart_tx_inst/r_Tx_Data [0]), 
            .I2(\uart_tx_inst/r_Bit_Index [2]), .O(n2827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8161.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8162 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .O(n2828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8162.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8163 (.I0(n2827), .I1(n2828), .I2(\uart_tx_inst/r_SM_Main [0]), 
            .I3(\uart_tx_inst/r_SM_Main [1]), .O(\uart_tx_inst/n634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40f */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(295)
    defparam LUT__8163.LUTMASK = 16'hf40f;
    EFX_LUT4 LUT__8164 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .O(\uart_tx_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(268)
    defparam LUT__8164.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8165 (.I0(\uart_tx_inst/LessThan_9/n18 ), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .I2(\uart_tx_inst/r_SM_Main [2]), .I3(\uart_tx_inst/r_SM_Main [0]), 
            .O(ceg_net28)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(211)
    defparam LUT__8165.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__8166 (.I0(\uart_tx_inst/r_SM_Main [1]), .I1(send), .O(n2829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8166.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8167 (.I0(\uart_tx_inst/r_SM_Main [0]), .I1(\uart_tx_inst/r_SM_Main [2]), 
            .I2(n2829), .O(\uart_tx_inst/n957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(51)
    defparam LUT__8167.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8168 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_Bit_Index [2]), .I3(\uart_tx_inst/r_SM_Main [1]), 
            .O(n2830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8168.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8169 (.I0(n2830), .I1(n2829), .I2(\uart_tx_inst/LessThan_9/n18 ), 
            .I3(\uart_tx_inst/r_SM_Main [0]), .O(\uart_tx_inst/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ce */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(295)
    defparam LUT__8169.LUTMASK = 16'hf0ce;
    EFX_LUT4 LUT__8170 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(n2826), .O(\uart_tx_inst/n716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8170.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8171 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .O(n2831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8171.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8172 (.I0(\uart_tx_inst/r_Clock_Count [2]), .I1(n2831), 
            .I2(n2826), .O(\uart_tx_inst/n719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8172.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8173 (.I0(\uart_tx_inst/r_Clock_Count [2]), .I1(n2831), 
            .I2(\uart_tx_inst/r_Clock_Count [3]), .I3(n2826), .O(\uart_tx_inst/n722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8173.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8174 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(\uart_tx_inst/r_Clock_Count [2]), .I3(\uart_tx_inst/r_Clock_Count [3]), 
            .O(n2832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8174.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8175 (.I0(\uart_tx_inst/r_Clock_Count [4]), .I1(n2832), 
            .I2(n2826), .O(\uart_tx_inst/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8175.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8176 (.I0(\uart_tx_inst/r_Clock_Count [4]), .I1(n2832), 
            .I2(\uart_tx_inst/r_Clock_Count [5]), .I3(n2826), .O(\uart_tx_inst/n728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8176.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8177 (.I0(n2824), .I1(n2832), .O(n2833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8177.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8178 (.I0(\uart_tx_inst/r_Clock_Count [6]), .I1(n2833), 
            .I2(n2826), .O(\uart_tx_inst/n731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8178.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8179 (.I0(\uart_tx_inst/r_Clock_Count [6]), .I1(n2833), 
            .O(n2834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8179.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8180 (.I0(\uart_tx_inst/r_Clock_Count [7]), .I1(n2834), 
            .I2(n2826), .O(\uart_tx_inst/n734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8180.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8181 (.I0(\uart_tx_inst/r_Clock_Count [7]), .I1(n2834), 
            .I2(\uart_tx_inst/r_Clock_Count [8]), .I3(n2826), .O(\uart_tx_inst/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(248)
    defparam LUT__8181.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__8182 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_SM_Main [1]), .O(\uart_tx_inst/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(268)
    defparam LUT__8182.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8183 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_Bit_Index [2]), .I3(\uart_tx_inst/r_SM_Main [1]), 
            .O(\uart_tx_inst/n814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(268)
    defparam LUT__8183.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__8184 (.I0(\uart_tx_inst/LessThan_9/n18 ), .I1(\uart_tx_inst/r_SM_Main [0]), 
            .I2(\uart_tx_inst/r_SM_Main [1]), .O(\uart_tx_inst/n709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(295)
    defparam LUT__8184.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__8185 (.I0(\uart_tx_inst/r_SM_Main [2]), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .I2(\uart_tx_inst/r_SM_Main [0]), .O(\uart_tx_inst/n945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(51)
    defparam LUT__8185.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__8186 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [5]), 
            .O(rx_data[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8186.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8187 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [6]), 
            .O(rx_data[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8187.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8188 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [7]), 
            .O(rx_data[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8188.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8191 (.I0(tx_2), .O(tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(296)
    defparam LUT__8191.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__8042 (.I0(\uart_rx_inst/r_Rx_Byte [0]), .I1(rx_ready), 
            .O(rx_data[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/add.v(179)
    defparam LUT__8042.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [0]), 
            .I1(1'b1), .CI(1'b0), .CO(n2835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4708)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_611fdb1c_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_611fdb1c_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_611fdb1c__5_5_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_611fdb1c_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_611fdb1c_0
// module not written out since it is a black box. 
//

