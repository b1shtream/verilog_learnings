
//
// Verific Verilog Description of module adder
//

module adder (clk, rx, tx, jtag_inst1_CAPTURE, jtag_inst1_DRCK, jtag_inst1_RESET, 
            jtag_inst1_RUNTEST, jtag_inst1_SEL, jtag_inst1_SHIFT, jtag_inst1_TCK, 
            jtag_inst1_TDI, jtag_inst1_TMS, jtag_inst1_UPDATE, jtag_inst1_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(2)
    input rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(3)
    output tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(4)
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire tx_2;
    wire [3:0]n25_2;
    wire [3:0]n30_2;
    wire [3:0]b;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(10)
    wire [3:0]sum;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(11)
    
    wire add_flag, send, carry;
    wire [3:0]a;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(10)
    
    wire \uart_rx_inst/r_Rx_Data , \uart_rx_inst/r_Rx_Data_R ;
    wire [8:0]\uart_rx_inst/r_Rx_Byte ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(74)
    wire [2:0]\uart_rx_inst/r_SM_Main ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(80)
    wire [31:0]\uart_rx_inst/r_Clock_Count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(72)
    
    wire rx_ready;
    wire [2:0]\uart_rx_inst/r_Bit_Index ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(73)
    wire [31:0]\uart_rx_inst/r_config_data ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(76)
    wire [31:0]\uart_tx_inst/r_Clock_Count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(195)
    wire [2:0]\uart_tx_inst/r_Bit_Index ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(196)
    wire [2:0]\uart_tx_inst/r_SM_Main ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(203)
    wire [31:0]\uart_tx_inst/r_config_data ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(200)
    wire [7:0]\uart_tx_inst/r_Tx_Data ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(197)
    
    wire \edb_top_inst/n1407 , \edb_top_inst/la0/la_run_trig ;
    wire [1:0]\edb_top_inst/la0/la_capture_pattern ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3438)
    wire [1:0]\edb_top_inst/la0/la_trig_pattern ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3426)
    
    wire \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig ;
    wire [255:0]\edb_top_inst/la0/la_trig_mask ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3433)
    wire [63:0]\edb_top_inst/la0/skip_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3428)
    wire [16:0]\edb_top_inst/la0/la_num_trigger ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3441)
    wire [4:0]\edb_top_inst/la0/la_window_depth ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3442)
    
    wire \edb_top_inst/la0/la_soft_reset_in ;
    wire [31:0]\edb_top_inst/la0/address_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3355)
    wire [3:0]\edb_top_inst/la0/opcode ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3354)
    wire [5:0]\edb_top_inst/la0/bit_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3356)
    wire [15:0]\edb_top_inst/la0/word_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3357)
    wire [63:0]\edb_top_inst/la0/data_out_shift_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3352)
    wire [3:0]\edb_top_inst/la0/module_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3412)
    
    wire \edb_top_inst/la0/la_resetn_p1 ;
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4190)
    
    wire \edb_top_inst/la0/la_resetn ;
    wire [0:0]\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4097)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4097)
    wire [2:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4190)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4206)
    wire [63:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4222)
    wire [8:0]\edb_top_inst/la0/cap_fifo_din_cu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3424)
    wire [8:0]\edb_top_inst/la0/cap_fifo_din_tu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3424)
    wire [12:0]\edb_top_inst/la0/internal_register_select ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3353)
    wire [16:0]\edb_top_inst/la0/la_trig_pos ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3421)
    wire [31:0]\edb_top_inst/la0/crc_data_out ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3408)
    
    wire \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ;
    wire [8:0]\edb_top_inst/la0/genblk4.cap_fifo_din_p1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4399)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5602)
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5602)
    
    wire \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/tu_trigger ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5819)
    
    wire \edb_top_inst/la0/ts_trigger ;
    wire [3:0]\edb_top_inst/la0/la_biu_inst/curr_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4903)
    
    wire \edb_top_inst/la0/la_biu_inst/run_trig_p2 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top_inst/la0/ts_resetn , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ;
    wire [63:0]\edb_top_inst/la0/data_from_biu ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3410)
    wire [1:0]\edb_top_inst/la0/la_biu_inst/axi_fsm_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4901)
    
    wire \edb_top_inst/la0/la_biu_inst/run_trig_p1 , \edb_top_inst/la0/biu_ready ;
    wire [31:0]\edb_top_inst/la0/la_biu_inst/addr_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4942)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5345)
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4606)
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4605)
    wire [16:0]\edb_top_inst/la0/la_sample_cnt ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3420)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4720)
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4935)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4596)
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4597)
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ;
    wire [3:0]\edb_top_inst/debug_hub_inst/module_id_reg ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(287)
    wire [81:0]\edb_top_inst/edb_user_dr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(33)
    wire [16:0]\edb_top_inst/la0/n1795 ;
    
    wire \edb_top_inst/la0/add_417/n2 ;
    wire [31:0]\edb_top_inst/la0/n1814 ;
    
    wire \edb_top_inst/la0/add_98/n2 ;
    wire [5:0]\edb_top_inst/la0/n1961 ;
    
    wire \edb_top_inst/la0/add_419/n2 ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/n73 ;
    
    wire \edb_top_inst/la0/trigger_skipper_n/add_19/n2 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n110 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ;
    wire [10:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 ;
    
    wire \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n124 , \edb_top_inst/la0/trigger_skipper_n/add_19/n122 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n120 , \edb_top_inst/la0/trigger_skipper_n/add_19/n118 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n116 , \edb_top_inst/la0/trigger_skipper_n/add_19/n114 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n112 , \edb_top_inst/la0/trigger_skipper_n/add_19/n110 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n108 , \edb_top_inst/la0/trigger_skipper_n/add_19/n106 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n104 , \edb_top_inst/la0/trigger_skipper_n/add_19/n102 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n100 , \edb_top_inst/la0/trigger_skipper_n/add_19/n98 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n96 , \edb_top_inst/la0/trigger_skipper_n/add_19/n94 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n92 , \edb_top_inst/la0/trigger_skipper_n/add_19/n90 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n88 , \edb_top_inst/la0/trigger_skipper_n/add_19/n86 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n84 , \edb_top_inst/la0/trigger_skipper_n/add_19/n82 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n80 , \edb_top_inst/la0/trigger_skipper_n/add_19/n78 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n76 , \edb_top_inst/la0/trigger_skipper_n/add_19/n74 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n72 , \edb_top_inst/la0/trigger_skipper_n/add_19/n70 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n68 , \edb_top_inst/la0/trigger_skipper_n/add_19/n66 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n64 , \edb_top_inst/la0/trigger_skipper_n/add_19/n62 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n60 , \edb_top_inst/la0/trigger_skipper_n/add_19/n58 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n56 , \edb_top_inst/la0/trigger_skipper_n/add_19/n54 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n52 , \edb_top_inst/la0/trigger_skipper_n/add_19/n50 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n48 , \edb_top_inst/la0/trigger_skipper_n/add_19/n46 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n44 , \edb_top_inst/la0/trigger_skipper_n/add_19/n42 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n40 , \edb_top_inst/la0/trigger_skipper_n/add_19/n38 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n36 , \edb_top_inst/la0/trigger_skipper_n/add_19/n34 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n32 , \edb_top_inst/la0/trigger_skipper_n/add_19/n30 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n28 , \edb_top_inst/la0/trigger_skipper_n/add_19/n26 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n24 , \edb_top_inst/la0/trigger_skipper_n/add_19/n22 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n20 , \edb_top_inst/la0/trigger_skipper_n/add_19/n18 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n16 , \edb_top_inst/la0/trigger_skipper_n/add_19/n14 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n12 , \edb_top_inst/la0/trigger_skipper_n/add_19/n10 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n8 , \edb_top_inst/la0/trigger_skipper_n/add_19/n6 , 
        \edb_top_inst/la0/trigger_skipper_n/add_19/n4 , \edb_top_inst/la0/add_419/n8 , 
        \edb_top_inst/la0/add_419/n6 , \edb_top_inst/la0/add_419/n4 , \edb_top_inst/la0/add_98/n48 , 
        \edb_top_inst/la0/add_98/n46 , \edb_top_inst/la0/add_98/n44 , \edb_top_inst/la0/add_98/n42 , 
        \edb_top_inst/la0/add_98/n40 , \edb_top_inst/la0/add_98/n38 , \edb_top_inst/la0/add_98/n36 , 
        \edb_top_inst/la0/add_98/n34 , \edb_top_inst/la0/add_98/n32 , \edb_top_inst/la0/add_98/n30 , 
        \edb_top_inst/la0/add_98/n28 , \edb_top_inst/la0/add_98/n26 , \edb_top_inst/la0/add_98/n24 , 
        \edb_top_inst/la0/add_98/n22 , \edb_top_inst/la0/add_98/n20 , \edb_top_inst/la0/add_98/n18 , 
        \edb_top_inst/la0/add_98/n16 , \edb_top_inst/la0/add_98/n14 , \edb_top_inst/la0/add_98/n12 , 
        \edb_top_inst/la0/add_98/n10 , \edb_top_inst/la0/add_98/n8 , \edb_top_inst/la0/add_98/n6 , 
        \edb_top_inst/la0/add_98/n4 , \edb_top_inst/la0/add_417/n16 , \edb_top_inst/la0/add_417/n14 , 
        \edb_top_inst/la0/add_417/n12 , \edb_top_inst/la0/add_417/n10 , 
        \edb_top_inst/la0/add_417/n8 , \edb_top_inst/la0/add_417/n6 , \edb_top_inst/la0/add_417/n4 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_dout ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4911)
    
    wire \edb_top_inst/n1408 , \edb_top_inst/n1409 , \edb_top_inst/n1410 , 
        \edb_top_inst/n1411 , \edb_top_inst/n1412 , \edb_top_inst/n1413 , 
        \edb_top_inst/n1414 , \edb_top_inst/n1415 , \edb_top_inst/n1416 , 
        \edb_top_inst/n1417 , \edb_top_inst/n1418 , \edb_top_inst/n1419 , 
        \edb_top_inst/n1420 , \edb_top_inst/n1421 , \edb_top_inst/n1422 , 
        \edb_top_inst/n1423 , \edb_top_inst/n1424 , \edb_top_inst/n1425 , 
        \edb_top_inst/n1426 , \edb_top_inst/n1427 , \edb_top_inst/n1428 , 
        \edb_top_inst/n1429 , \edb_top_inst/n1430 , \edb_top_inst/n1431 , 
        \edb_top_inst/n1432 , \edb_top_inst/n1433 , \edb_top_inst/n1434 , 
        \edb_top_inst/n1435 , \edb_top_inst/n1436 , \edb_top_inst/n1437 , 
        \edb_top_inst/n1438 , \edb_top_inst/n1439 , \edb_top_inst/n1440 , 
        \edb_top_inst/n1441 , \edb_top_inst/n1442 , \edb_top_inst/n1443 , 
        \edb_top_inst/n1444 , \edb_top_inst/n1445 , \edb_top_inst/n1446 , 
        \edb_top_inst/n1447 , \edb_top_inst/n1448 , \edb_top_inst/n1449 , 
        \edb_top_inst/n1450 , \edb_top_inst/n1451 , \edb_top_inst/la0/n999 , 
        \edb_top_inst/n1452 , \edb_top_inst/n1453 , \edb_top_inst/n1454 , 
        \edb_top_inst/n1455 , \edb_top_inst/n1456 , \edb_top_inst/la0/regsel_ld_en , 
        \edb_top_inst/n1457 , \edb_top_inst/n1458 , \edb_top_inst/n1459 , 
        \edb_top_inst/la0/n971 , \edb_top_inst/ceg_net2 , \edb_top_inst/la0/n1000 , 
        \edb_top_inst/la0/n1001 , \edb_top_inst/la0/n1055 , \edb_top_inst/n1460 , 
        \edb_top_inst/la0/n1572 , \edb_top_inst/la0/n1705 , \edb_top_inst/n1461 , 
        \edb_top_inst/n1462 , \edb_top_inst/la0/n1757 , \edb_top_inst/n1463 , 
        \edb_top_inst/n1464 , \edb_top_inst/n1465 , \edb_top_inst/n1466 , 
        \edb_top_inst/n1467 ;
    wire [31:0]\edb_top_inst/la0/data_to_addr_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3402)
    
    wire \edb_top_inst/la0/op_reg_en , \edb_top_inst/n1468 , \edb_top_inst/n1469 , 
        \edb_top_inst/n1470 , \edb_top_inst/la0/n595 , \edb_top_inst/la0/n596 , 
        \edb_top_inst/n1471 , \edb_top_inst/n1472 , \edb_top_inst/n1473 , 
        \edb_top_inst/la0/n593 , \edb_top_inst/n1474 , \edb_top_inst/n1475 , 
        \edb_top_inst/n1476 , \edb_top_inst/n1477 , \edb_top_inst/n1478 , 
        \edb_top_inst/n1479 , \edb_top_inst/n1480 , \edb_top_inst/n1481 , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/n1482 , \edb_top_inst/n1483 , 
        \edb_top_inst/n1484 ;
    wire [5:0]\edb_top_inst/la0/n1975 ;
    
    wire \edb_top_inst/n1485 , \edb_top_inst/n1486 , \edb_top_inst/n1487 , 
        \edb_top_inst/n1488 , \edb_top_inst/n1489 ;
    wire [3:0]\edb_top_inst/la0/module_next_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3412)
    
    wire \edb_top_inst/n1490 , \edb_top_inst/ceg_net5 ;
    wire [15:0]\edb_top_inst/la0/data_to_word_counter ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3405)
    
    wire \edb_top_inst/n1491 , \edb_top_inst/la0/word_ct_en , \edb_top_inst/n1492 , 
        \edb_top_inst/n1493 , \edb_top_inst/n1494 , \edb_top_inst/n1495 , 
        \edb_top_inst/n1496 , \edb_top_inst/n1497 , \edb_top_inst/n1498 , 
        \edb_top_inst/n1499 , \edb_top_inst/n1500 , \edb_top_inst/n1501 , 
        \edb_top_inst/n1502 , \edb_top_inst/n1503 , \edb_top_inst/n1504 , 
        \edb_top_inst/n1505 , \edb_top_inst/n1506 , \edb_top_inst/n1507 , 
        \edb_top_inst/n1508 ;
    wire [63:0]\edb_top_inst/la0/n2194 ;
    
    wire \edb_top_inst/n1509 , \edb_top_inst/ceg_net8 , \edb_top_inst/la0/n2545 , 
        \edb_top_inst/la0/n2558 , \edb_top_inst/n1510 , \edb_top_inst/la0/n3447 , 
        \edb_top_inst/la0/n3462 , \edb_top_inst/la0/n3660 , \edb_top_inst/n1511 , 
        \edb_top_inst/n1512 , \edb_top_inst/n1513 , \edb_top_inst/n1514 , 
        \edb_top_inst/n1515 , \edb_top_inst/n1516 , \edb_top_inst/n1517 , 
        \edb_top_inst/n1518 , \edb_top_inst/n1519 , \edb_top_inst/n1520 , 
        \edb_top_inst/n1528 , \edb_top_inst/n1529 , \edb_top_inst/n1530 , 
        \edb_top_inst/n1531 , \edb_top_inst/n1532 , \edb_top_inst/n1533 , 
        \edb_top_inst/n1534 , \edb_top_inst/n1535 , \edb_top_inst/n1536 , 
        \edb_top_inst/n1537 , \edb_top_inst/n1538 , \edb_top_inst/n1539 , 
        \edb_top_inst/n1540 , \edb_top_inst/n1541 , \edb_top_inst/n1542 , 
        \edb_top_inst/n1544 , \edb_top_inst/n1545 , \edb_top_inst/n1546 , 
        \edb_top_inst/n1547 , \edb_top_inst/n1548 , \edb_top_inst/n1549 , 
        \edb_top_inst/n1550 , \edb_top_inst/n1551 , \edb_top_inst/n1552 , 
        \edb_top_inst/n1553 , \edb_top_inst/n1554 , \edb_top_inst/n1555 , 
        \edb_top_inst/n1556 , \edb_top_inst/n1557 , \edb_top_inst/n1558 , 
        \edb_top_inst/n1559 , \edb_top_inst/n1560 , \edb_top_inst/n1561 , 
        \edb_top_inst/n1562 , \edb_top_inst/n1563 , \edb_top_inst/n1564 , 
        \edb_top_inst/n1565 , \edb_top_inst/n1566 , \edb_top_inst/n1567 , 
        \edb_top_inst/n1568 , \edb_top_inst/n1569 , \edb_top_inst/n1570 , 
        \edb_top_inst/n1571 , \edb_top_inst/n1572 , \edb_top_inst/n1573 , 
        \edb_top_inst/n1574 , \edb_top_inst/n1575 , \edb_top_inst/n1576 , 
        \edb_top_inst/n1577 , \edb_top_inst/n1578 , \edb_top_inst/n1579 , 
        \edb_top_inst/n1580 , \edb_top_inst/n1581 , \edb_top_inst/n1582 , 
        \edb_top_inst/n1583 , \edb_top_inst/n1584 , \edb_top_inst/n1585 , 
        \edb_top_inst/n1586 , \edb_top_inst/n1587 , \edb_top_inst/n1588 , 
        \edb_top_inst/n1589 , \edb_top_inst/n1590 , \edb_top_inst/n1591 , 
        \edb_top_inst/n1592 , \edb_top_inst/n1593 , \edb_top_inst/n1594 , 
        \edb_top_inst/n1595 , \edb_top_inst/n1596 , \edb_top_inst/n1597 , 
        \edb_top_inst/n1598 , \edb_top_inst/n1599 , \edb_top_inst/n1600 , 
        \edb_top_inst/n1601 , \edb_top_inst/n1602 , \edb_top_inst/n1604 , 
        \edb_top_inst/n1605 , \edb_top_inst/n1606 , \edb_top_inst/n1607 , 
        \edb_top_inst/n1608 , \edb_top_inst/n1609 , \edb_top_inst/n1610 , 
        \edb_top_inst/n1611 , \edb_top_inst/n1612 , \edb_top_inst/n1613 , 
        \edb_top_inst/n1614 , \edb_top_inst/n1615 , \edb_top_inst/n1616 , 
        \edb_top_inst/n1617 , \edb_top_inst/n1618 , \edb_top_inst/n1619 , 
        \edb_top_inst/n1620 , \edb_top_inst/n1621 , \edb_top_inst/n1622 , 
        \edb_top_inst/n1623 , \edb_top_inst/n1624 , \edb_top_inst/n1625 , 
        \edb_top_inst/n1626 , \edb_top_inst/n1627 , \edb_top_inst/n1628 , 
        \edb_top_inst/n1629 , \edb_top_inst/n1630 , \edb_top_inst/n1631 , 
        \edb_top_inst/n1632 , \edb_top_inst/n1633 , \edb_top_inst/n1634 , 
        \edb_top_inst/n1635 , \edb_top_inst/n1636 , \edb_top_inst/n1637 , 
        \edb_top_inst/n1638 , \edb_top_inst/n1639 , \edb_top_inst/n1640 , 
        \edb_top_inst/n1641 , \edb_top_inst/n1642 , \edb_top_inst/n1643 , 
        \edb_top_inst/n1644 , \edb_top_inst/n1645 , \edb_top_inst/n1646 , 
        \edb_top_inst/n1647 , \edb_top_inst/n1648 , \edb_top_inst/n1649 , 
        \edb_top_inst/n1651 , \edb_top_inst/n1652 , \edb_top_inst/n1653 , 
        \edb_top_inst/n1654 , \edb_top_inst/n1655 , \edb_top_inst/n1656 , 
        \edb_top_inst/n1657 , \edb_top_inst/n1658 , \edb_top_inst/n1659 , 
        \edb_top_inst/n1660 , \edb_top_inst/n1661 , \edb_top_inst/n1662 , 
        \edb_top_inst/n1663 , \edb_top_inst/n1664 , \edb_top_inst/n1665 , 
        \edb_top_inst/n1666 , \edb_top_inst/n1667 , \edb_top_inst/n1668 , 
        \edb_top_inst/n1669 , \edb_top_inst/n1670 , \edb_top_inst/n1671 , 
        \edb_top_inst/n1672 , \edb_top_inst/n1673 , \edb_top_inst/n1674 , 
        \edb_top_inst/n1675 , \edb_top_inst/n1676 , \edb_top_inst/n1677 , 
        \edb_top_inst/n1678 , \edb_top_inst/n1679 , \edb_top_inst/n1680 , 
        \edb_top_inst/n1681 , \edb_top_inst/n1682 , \edb_top_inst/n1683 , 
        \edb_top_inst/n1684 , \edb_top_inst/n1685 , \edb_top_inst/n1686 , 
        \edb_top_inst/n1687 , \edb_top_inst/n1688 ;
    wire [31:0]\edb_top_inst/la0/axi_crc_i/n118 ;
    
    wire \edb_top_inst/n1689 , \edb_top_inst/ceg_net11 , \edb_top_inst/n1690 , 
        \edb_top_inst/n1691 , \edb_top_inst/n1692 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n1693 , \edb_top_inst/n1694 , \edb_top_inst/n1695 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 ;
    wire [7:0]\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 ;
    
    wire \edb_top_inst/n1696 , \edb_top_inst/n1697 , \edb_top_inst/n1698 , 
        \edb_top_inst/n1699 , \edb_top_inst/n1700 , \edb_top_inst/n1701 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/n1702 , 
        \edb_top_inst/n1703 , \edb_top_inst/n1704 , \edb_top_inst/n1705 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/n1706 , \edb_top_inst/n1707 , \edb_top_inst/n1708 , 
        \edb_top_inst/n1709 , \edb_top_inst/n1710 , \edb_top_inst/n1711 , 
        \edb_top_inst/n1712 , \edb_top_inst/n1713 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/n1714 , \edb_top_inst/n1715 , \edb_top_inst/n1716 , 
        \edb_top_inst/la0/trigger_tu/n29 , \edb_top_inst/n1717 , \edb_top_inst/n1718 , 
        \edb_top_inst/n1719 , \edb_top_inst/n1720 , \edb_top_inst/n1721 , 
        \edb_top_inst/n1722 , \edb_top_inst/n1723 , \edb_top_inst/n1724 , 
        \edb_top_inst/n1725 , \edb_top_inst/n1726 , \edb_top_inst/n1727 , 
        \edb_top_inst/n1728 , \edb_top_inst/n1729 , \edb_top_inst/n1730 , 
        \edb_top_inst/n1731 , \edb_top_inst/n1732 , \edb_top_inst/n1733 , 
        \edb_top_inst/n1734 , \edb_top_inst/n1735 , \edb_top_inst/n1736 , 
        \edb_top_inst/n1737 , \edb_top_inst/n1738 , \edb_top_inst/n1739 , 
        \edb_top_inst/n1740 , \edb_top_inst/n1741 , \edb_top_inst/n1742 , 
        \edb_top_inst/n1743 , \edb_top_inst/n1744 , \edb_top_inst/n1745 , 
        \edb_top_inst/n1746 , \edb_top_inst/n1747 , \edb_top_inst/n1748 , 
        \edb_top_inst/n1749 , \edb_top_inst/n1750 , \edb_top_inst/n1751 , 
        \edb_top_inst/n1752 , \edb_top_inst/n1753 , \edb_top_inst/n1754 , 
        \edb_top_inst/n1755 , \edb_top_inst/n1756 , \edb_top_inst/n1757 , 
        \edb_top_inst/n1758 , \edb_top_inst/n1759 , \edb_top_inst/n1760 , 
        \edb_top_inst/n1761 , \edb_top_inst/n1762 , \edb_top_inst/n1763 , 
        \edb_top_inst/n1764 , \edb_top_inst/n1765 , \edb_top_inst/n1766 , 
        \edb_top_inst/n1767 , \edb_top_inst/n1768 , \edb_top_inst/n1769 , 
        \edb_top_inst/n1770 , \edb_top_inst/n1771 , \edb_top_inst/n1772 , 
        \edb_top_inst/n1773 , \edb_top_inst/n1774 , \edb_top_inst/n1775 , 
        \edb_top_inst/n1776 , \edb_top_inst/n1777 , \edb_top_inst/n1778 , 
        \edb_top_inst/n1779 , \edb_top_inst/n1780 , \edb_top_inst/n1781 , 
        \edb_top_inst/n1782 , \edb_top_inst/n1783 , \edb_top_inst/n1784 , 
        \edb_top_inst/n1785 , \edb_top_inst/n1786 , \edb_top_inst/n1787 , 
        \edb_top_inst/n1788 , \edb_top_inst/n1789 , \edb_top_inst/n1790 , 
        \edb_top_inst/n1791 , \edb_top_inst/n1792 , \edb_top_inst/n1793 , 
        \edb_top_inst/n1794 , \edb_top_inst/n1795 , \edb_top_inst/n1796 , 
        \edb_top_inst/n1797 , \edb_top_inst/n1798 , \edb_top_inst/n1799 , 
        \edb_top_inst/n1800 , \edb_top_inst/n1801 , \edb_top_inst/n1802 , 
        \edb_top_inst/n1803 , \edb_top_inst/n1804 , \edb_top_inst/n1805 , 
        \edb_top_inst/n1806 , \edb_top_inst/n1807 , \edb_top_inst/n1808 , 
        \edb_top_inst/n1809 , \edb_top_inst/n1810 , \edb_top_inst/n1811 , 
        \edb_top_inst/n1812 , \edb_top_inst/n1813 , \edb_top_inst/n1814 , 
        \edb_top_inst/n1815 , \edb_top_inst/n1816 , \edb_top_inst/n1817 , 
        \edb_top_inst/n1818 , \edb_top_inst/n1819 , \edb_top_inst/n1820 , 
        \edb_top_inst/n1821 , \edb_top_inst/n1822 , \edb_top_inst/n1823 , 
        \edb_top_inst/n1824 , \edb_top_inst/n1825 , \edb_top_inst/n1826 , 
        \edb_top_inst/n1827 , \edb_top_inst/n1828 , \edb_top_inst/n1829 , 
        \edb_top_inst/n1830 , \edb_top_inst/n1831 , \edb_top_inst/n1832 , 
        \edb_top_inst/n1833 , \edb_top_inst/n1834 , \edb_top_inst/n1835 , 
        \edb_top_inst/n1836 , \edb_top_inst/n1837 , \edb_top_inst/n1838 , 
        \edb_top_inst/n1839 , \edb_top_inst/n1840 , \edb_top_inst/n1841 , 
        \edb_top_inst/n1842 , \edb_top_inst/n1843 , \edb_top_inst/n1844 , 
        \edb_top_inst/n1845 , \edb_top_inst/n1846 , \edb_top_inst/n1847 , 
        \edb_top_inst/n1848 , \edb_top_inst/n1849 , \edb_top_inst/n1850 , 
        \edb_top_inst/n1851 , \edb_top_inst/n1852 , \edb_top_inst/n1853 , 
        \edb_top_inst/n1854 , \edb_top_inst/n1855 , \edb_top_inst/n1856 , 
        \edb_top_inst/n1857 , \edb_top_inst/n1858 , \edb_top_inst/n1859 , 
        \edb_top_inst/n1860 , \edb_top_inst/n1861 , \edb_top_inst/n1862 , 
        \edb_top_inst/n1863 , \edb_top_inst/n1864 , \edb_top_inst/n1865 , 
        \edb_top_inst/n1866 , \edb_top_inst/n1867 , \edb_top_inst/n1868 , 
        \edb_top_inst/n1869 , \edb_top_inst/n1870 , \edb_top_inst/n1871 , 
        \edb_top_inst/n1872 , \edb_top_inst/n1873 , \edb_top_inst/n1874 , 
        \edb_top_inst/n1875 , \edb_top_inst/n1876 , \edb_top_inst/n1877 ;
    wire [63:0]\edb_top_inst/la0/trigger_skipper_n/n138 ;
    
    wire \edb_top_inst/la0/trigger_skipper_n/n468 , \edb_top_inst/n1878 , 
        \edb_top_inst/n1879 , \edb_top_inst/n1880 , \edb_top_inst/n1881 , 
        \edb_top_inst/n1882 , \edb_top_inst/n1883 , \edb_top_inst/n1884 , 
        \edb_top_inst/n1885 , \edb_top_inst/n1886 , \edb_top_inst/n1887 , 
        \edb_top_inst/n1888 , \edb_top_inst/n1889 , \edb_top_inst/n1890 , 
        \edb_top_inst/n1891 , \edb_top_inst/n1892 , \edb_top_inst/n1893 , 
        \edb_top_inst/n1894 , \edb_top_inst/n1895 , \edb_top_inst/n1896 , 
        \edb_top_inst/n1897 , \edb_top_inst/n1898 , \edb_top_inst/n1899 , 
        \edb_top_inst/n1900 , \edb_top_inst/n1901 , \edb_top_inst/n1902 , 
        \edb_top_inst/n1903 , \edb_top_inst/n1904 , \edb_top_inst/n1905 , 
        \edb_top_inst/n1906 , \edb_top_inst/n1907 , \edb_top_inst/n1908 , 
        \edb_top_inst/n1909 , \edb_top_inst/n1910 , \edb_top_inst/n1911 , 
        \edb_top_inst/n1912 , \edb_top_inst/n1913 , \edb_top_inst/n1914 , 
        \edb_top_inst/n1915 , \edb_top_inst/n1916 , \edb_top_inst/n1917 , 
        \edb_top_inst/n1918 , \edb_top_inst/n1919 , \edb_top_inst/n1920 , 
        \edb_top_inst/n1921 , \edb_top_inst/n1922 , \edb_top_inst/n1923 , 
        \edb_top_inst/n1924 , \edb_top_inst/n1925 , \edb_top_inst/n1926 , 
        \edb_top_inst/n1927 , \edb_top_inst/n1928 , \edb_top_inst/n1929 , 
        \edb_top_inst/n1930 , \edb_top_inst/n1931 , \edb_top_inst/n1932 , 
        \edb_top_inst/n1933 , \edb_top_inst/n1934 , \edb_top_inst/n1935 , 
        \edb_top_inst/n1936 , \edb_top_inst/n1937 , \edb_top_inst/n1938 , 
        \edb_top_inst/n1939 , \edb_top_inst/n1940 , \edb_top_inst/n1941 , 
        \edb_top_inst/n1942 , \edb_top_inst/n1943 , \edb_top_inst/n1944 , 
        \edb_top_inst/n1945 , \edb_top_inst/n1946 , \edb_top_inst/n1947 , 
        \edb_top_inst/n1948 , \edb_top_inst/n1949 , \edb_top_inst/n1950 , 
        \edb_top_inst/n1951 , \edb_top_inst/n1952 , \edb_top_inst/n1953 , 
        \edb_top_inst/n1954 , \edb_top_inst/n1955 , \edb_top_inst/n1956 , 
        \edb_top_inst/n1957 , \edb_top_inst/n1958 , \edb_top_inst/n1959 , 
        \edb_top_inst/n1960 , \edb_top_inst/n1961 , \edb_top_inst/n1962 , 
        \edb_top_inst/n1963 , \edb_top_inst/n1964 , \edb_top_inst/n1965 , 
        \edb_top_inst/n1966 , \edb_top_inst/n1967 , \edb_top_inst/n1968 , 
        \edb_top_inst/n1969 , \edb_top_inst/n1970 , \edb_top_inst/n1971 , 
        \edb_top_inst/n1972 , \edb_top_inst/n1973 , \edb_top_inst/n1974 , 
        \edb_top_inst/n1975 , \edb_top_inst/n1976 , \edb_top_inst/n1977 , 
        \edb_top_inst/n1978 , \edb_top_inst/n1979 , \edb_top_inst/n1980 , 
        \edb_top_inst/n1981 , \edb_top_inst/n1982 , \edb_top_inst/n1983 , 
        \edb_top_inst/n1984 , \edb_top_inst/n1985 , \edb_top_inst/n1986 , 
        \edb_top_inst/n1987 , \edb_top_inst/n1988 , \edb_top_inst/n1989 , 
        \edb_top_inst/n1990 , \edb_top_inst/n1991 , \edb_top_inst/n1992 , 
        \edb_top_inst/n1993 , \edb_top_inst/n1994 , \edb_top_inst/n1995 , 
        \edb_top_inst/n1996 , \edb_top_inst/n1997 , \edb_top_inst/n1998 ;
    wire [3:0]\edb_top_inst/la0/la_biu_inst/next_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4903)
    
    wire \edb_top_inst/la0/la_biu_inst/n63 , \edb_top_inst/la0/la_biu_inst/n335 , 
        \edb_top_inst/la0/la_biu_inst/n1248 , \edb_top_inst/la0/la_biu_inst/n1249 , 
        \edb_top_inst/la0/la_biu_inst/n1832 , \edb_top_inst/n1999 , \edb_top_inst/n2000 , 
        \edb_top_inst/la0/la_biu_inst/n1214 , \edb_top_inst/la0/n5970 , 
        \edb_top_inst/n2001 , \edb_top_inst/n2002 , \edb_top_inst/n2003 , 
        \edb_top_inst/n2004 , \edb_top_inst/n2005 , \edb_top_inst/n2006 , 
        \edb_top_inst/n2007 , \edb_top_inst/n2008 , \edb_top_inst/n2009 , 
        \edb_top_inst/n2010 , \edb_top_inst/n2011 , \edb_top_inst/n2012 , 
        \edb_top_inst/n2013 , \edb_top_inst/n2014 , \edb_top_inst/ceg_net18 ;
    wire [1:0]\edb_top_inst/la0/la_biu_inst/next_fsm_state ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4901)
    
    wire \edb_top_inst/ceg_net24 , \edb_top_inst/n2015 , \edb_top_inst/la0/la_biu_inst/n1839 , 
        \edb_top_inst/la0/la_biu_inst/fifo_push , \edb_top_inst/n2016 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , \edb_top_inst/la0/la_biu_inst/fifo_rstn , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 , \edb_top_inst/~ceg_net27 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n576 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , \edb_top_inst/n2017 , 
        \edb_top_inst/n2018 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4533)
    
    wire \edb_top_inst/n2019 , \edb_top_inst/n2020 , \edb_top_inst/n2021 , 
        \edb_top_inst/n2022 , \edb_top_inst/n2023 , \edb_top_inst/n2024 , 
        \edb_top_inst/n2025 , \edb_top_inst/n2026 , \edb_top_inst/n2027 , 
        \edb_top_inst/n2028 , \edb_top_inst/n2029 , \edb_top_inst/n2030 , 
        \edb_top_inst/n2031 , \edb_top_inst/n2032 , \edb_top_inst/n2033 , 
        \edb_top_inst/n2034 , \edb_top_inst/n2035 , \edb_top_inst/n2036 , 
        \edb_top_inst/n2037 , \edb_top_inst/n2038 , \edb_top_inst/n2039 , 
        \edb_top_inst/n2040 , \edb_top_inst/n2041 , \edb_top_inst/n2042 , 
        \edb_top_inst/n2043 , \edb_top_inst/n2044 , \edb_top_inst/n2045 , 
        \edb_top_inst/n2046 , \edb_top_inst/n2047 , \edb_top_inst/n2048 , 
        \edb_top_inst/n2049 , \edb_top_inst/n2050 ;
    wire [9:0]\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4533)
    
    wire \edb_top_inst/la0/n594 , \edb_top_inst/n2051 , \edb_top_inst/debug_hub_inst/n266 , 
        \edb_top_inst/debug_hub_inst/n95 , \edb_top_inst/n1406 , n2336;
    wire [7:0]rx_data;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(7)
    
    wire \uart_rx_inst/n1220 , \uart_rx_inst/n1145 , \uart_rx_inst/n1148 , 
        ceg_net14, \uart_rx_inst/n337 , ceg_net32, \uart_rx_inst/n1152 , 
        ceg_net26, \uart_rx_inst/n1199 , \uart_rx_inst/n1202 , \uart_rx_inst/n1205 , 
        \uart_rx_inst/n1208 , \uart_rx_inst/n1211 , \uart_rx_inst/n1214 , 
        \uart_rx_inst/n1217 , \uart_rx_inst/n826 , \uart_rx_inst/n151 , 
        \uart_rx_inst/n1180 , \uart_rx_inst/n833 , \uart_rx_inst/n836 , 
        \uart_rx_inst/n839 , \uart_rx_inst/n842 , \uart_rx_inst/n845 , 
        \uart_rx_inst/n848 , \uart_rx_inst/n851 , \uart_rx_inst/n854 , 
        \uart_rx_inst/n857 , \uart_rx_inst/n860 , \uart_rx_inst/n863 , 
        \uart_rx_inst/n866 , \uart_rx_inst/n869 , \uart_rx_inst/n872 , 
        \uart_rx_inst/n875 , \uart_rx_inst/n878 , \uart_rx_inst/n881 , 
        \uart_rx_inst/n884 , \uart_rx_inst/n887 , \uart_rx_inst/n890 , 
        \uart_rx_inst/n893 , \uart_rx_inst/n896 , \uart_rx_inst/n899 , 
        \uart_rx_inst/n902 , \uart_rx_inst/n905 , \uart_rx_inst/n908 , 
        \uart_rx_inst/n911 , \uart_rx_inst/n914 , \uart_rx_inst/n917 , 
        \uart_rx_inst/n920 , \uart_rx_inst/n923 , \uart_rx_inst/n927 , 
        \uart_rx_inst/n931 , \uart_rx_inst/n1161 ;
    wire [3:0]n25;
    
    wire \uart_tx_inst/n1116 , \uart_tx_inst/n733 , \uart_tx_inst/n1120 , 
        ceg_net28, \uart_tx_inst/n1112 , \uart_tx_inst/n786 , \uart_tx_inst/n789 , 
        \uart_tx_inst/n792 , \uart_tx_inst/n795 , \uart_tx_inst/n798 , 
        \uart_tx_inst/n801 , \uart_tx_inst/n804 , \uart_tx_inst/n807 , 
        \uart_tx_inst/n810 , \uart_tx_inst/n813 , \uart_tx_inst/n816 , 
        \uart_tx_inst/n819 , \uart_tx_inst/n822 , \uart_tx_inst/n825 , 
        \uart_tx_inst/n828 , \uart_tx_inst/n831 , \uart_tx_inst/n834 , 
        \uart_tx_inst/n837 , \uart_tx_inst/n840 , \uart_tx_inst/n843 , 
        \uart_tx_inst/n846 , \uart_tx_inst/n849 , \uart_tx_inst/n852 , 
        \uart_tx_inst/n855 , \uart_tx_inst/n858 , \uart_tx_inst/n861 , 
        \uart_tx_inst/n864 , \uart_tx_inst/n867 , \uart_tx_inst/n870 , 
        \uart_tx_inst/n873 , \uart_tx_inst/n876 , \uart_tx_inst/n880 , 
        \uart_tx_inst/n884 , \uart_tx_inst/n1032 , \uart_tx_inst/n1224 , 
        \uart_tx_inst/n779 , \uart_tx_inst/n50 , \uart_tx_inst/n1206 , 
        \jtag_inst1_TCK~O , \clk~O , n2337, n2195, n2196, n2197, 
        n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
        n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
        n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, 
        n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
        n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
        n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
        n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
        n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, 
        n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
        n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
        n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
        n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
        n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
        n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
        n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, 
        n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
        n2334, n2335;
    
    EFX_LUT4 LUT__6230 (.I0(b[0]), .I1(a[0]), .O(n25_2[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(35)
    defparam LUT__6230.LUTMASK = 16'h6666;
    EFX_FF \b[0]~FF  (.D(rx_data[0]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \b[0]~FF .CLK_POLARITY = 1'b1;
    defparam \b[0]~FF .CE_POLARITY = 1'b1;
    defparam \b[0]~FF .SR_POLARITY = 1'b1;
    defparam \b[0]~FF .D_POLARITY = 1'b1;
    defparam \b[0]~FF .SR_SYNC = 1'b1;
    defparam \b[0]~FF .SR_VALUE = 1'b0;
    defparam \b[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \sum[0]~FF  (.D(n25_2[0]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(sum[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \sum[0]~FF .CLK_POLARITY = 1'b1;
    defparam \sum[0]~FF .CE_POLARITY = 1'b1;
    defparam \sum[0]~FF .SR_POLARITY = 1'b1;
    defparam \sum[0]~FF .D_POLARITY = 1'b1;
    defparam \sum[0]~FF .SR_SYNC = 1'b1;
    defparam \sum[0]~FF .SR_VALUE = 1'b0;
    defparam \sum[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \add_flag~FF  (.D(1'b1), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(add_flag)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \add_flag~FF .CLK_POLARITY = 1'b1;
    defparam \add_flag~FF .CE_POLARITY = 1'b1;
    defparam \add_flag~FF .SR_POLARITY = 1'b1;
    defparam \add_flag~FF .D_POLARITY = 1'b1;
    defparam \add_flag~FF .SR_SYNC = 1'b1;
    defparam \add_flag~FF .SR_VALUE = 1'b0;
    defparam \add_flag~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \send~FF  (.D(1'b1), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(send)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \send~FF .CLK_POLARITY = 1'b1;
    defparam \send~FF .CE_POLARITY = 1'b1;
    defparam \send~FF .SR_POLARITY = 1'b1;
    defparam \send~FF .D_POLARITY = 1'b1;
    defparam \send~FF .SR_SYNC = 1'b1;
    defparam \send~FF .SR_VALUE = 1'b0;
    defparam \send~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \carry~FF  (.D(n30_2[0]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(carry)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \carry~FF .CLK_POLARITY = 1'b1;
    defparam \carry~FF .CE_POLARITY = 1'b1;
    defparam \carry~FF .SR_POLARITY = 1'b1;
    defparam \carry~FF .D_POLARITY = 1'b1;
    defparam \carry~FF .SR_SYNC = 1'b1;
    defparam \carry~FF .SR_VALUE = 1'b0;
    defparam \carry~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[0]~FF  (.D(rx_data[4]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \a[0]~FF .CLK_POLARITY = 1'b1;
    defparam \a[0]~FF .CE_POLARITY = 1'b1;
    defparam \a[0]~FF .SR_POLARITY = 1'b1;
    defparam \a[0]~FF .D_POLARITY = 1'b1;
    defparam \a[0]~FF .SR_SYNC = 1'b1;
    defparam \a[0]~FF .SR_VALUE = 1'b0;
    defparam \a[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Data~FF  (.D(\uart_rx_inst/r_Rx_Data_R ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(94)
    defparam \uart_rx_inst/r_Rx_Data~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Data_R~FF  (.D(rx), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Data_R )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Data_R~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Data_R~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[0]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1220 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[0]~FF  (.D(\uart_rx_inst/n1145 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/r_SM_Main [2]), .Q(\uart_rx_inst/r_SM_Main [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[0]~FF  (.D(\uart_rx_inst/n1148 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_ready~FF  (.D(\uart_rx_inst/n337 ), .CE(ceg_net32), .CLK(\clk~O ), 
           .SR(1'b0), .Q(rx_ready)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \rx_ready~FF .CLK_POLARITY = 1'b1;
    defparam \rx_ready~FF .CE_POLARITY = 1'b0;
    defparam \rx_ready~FF .SR_POLARITY = 1'b1;
    defparam \rx_ready~FF .D_POLARITY = 1'b1;
    defparam \rx_ready~FF .SR_SYNC = 1'b1;
    defparam \rx_ready~FF .SR_VALUE = 1'b0;
    defparam \rx_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[0]~FF  (.D(\uart_rx_inst/n1152 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[1]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1199 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[2]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[3]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1205 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[4]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1208 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[5]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1211 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[6]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1214 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Rx_Byte[7]~FF  (.D(\uart_rx_inst/r_Rx_Data ), .CE(\uart_rx_inst/n1217 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Rx_Byte [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Rx_Byte[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[1]~FF  (.D(\uart_rx_inst/n826 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/r_SM_Main [2]), .Q(\uart_rx_inst/r_SM_Main [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_SM_Main[2]~FF  (.D(\uart_rx_inst/n151 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_rx_inst/n1180 ), .Q(\uart_rx_inst/r_SM_Main [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[1]~FF  (.D(\uart_rx_inst/n833 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[2]~FF  (.D(\uart_rx_inst/n836 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[3]~FF  (.D(\uart_rx_inst/n839 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[4]~FF  (.D(\uart_rx_inst/n842 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[5]~FF  (.D(\uart_rx_inst/n845 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[6]~FF  (.D(\uart_rx_inst/n848 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[7]~FF  (.D(\uart_rx_inst/n851 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[8]~FF  (.D(\uart_rx_inst/n854 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[9]~FF  (.D(\uart_rx_inst/n857 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[10]~FF  (.D(\uart_rx_inst/n860 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[11]~FF  (.D(\uart_rx_inst/n863 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[12]~FF  (.D(\uart_rx_inst/n866 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[13]~FF  (.D(\uart_rx_inst/n869 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[14]~FF  (.D(\uart_rx_inst/n872 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[15]~FF  (.D(\uart_rx_inst/n875 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[16]~FF  (.D(\uart_rx_inst/n878 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[17]~FF  (.D(\uart_rx_inst/n881 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[18]~FF  (.D(\uart_rx_inst/n884 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[19]~FF  (.D(\uart_rx_inst/n887 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[20]~FF  (.D(\uart_rx_inst/n890 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[21]~FF  (.D(\uart_rx_inst/n893 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[22]~FF  (.D(\uart_rx_inst/n896 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[23]~FF  (.D(\uart_rx_inst/n899 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[24]~FF  (.D(\uart_rx_inst/n902 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[25]~FF  (.D(\uart_rx_inst/n905 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[26]~FF  (.D(\uart_rx_inst/n908 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[27]~FF  (.D(\uart_rx_inst/n911 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[28]~FF  (.D(\uart_rx_inst/n914 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[29]~FF  (.D(\uart_rx_inst/n917 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[30]~FF  (.D(\uart_rx_inst/n920 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Clock_Count[31]~FF  (.D(\uart_rx_inst/n923 ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Clock_Count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Clock_Count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[1]~FF  (.D(\uart_rx_inst/n927 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_Bit_Index[2]~FF  (.D(\uart_rx_inst/n931 ), .CE(ceg_net26), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_Bit_Index [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx_inst/r_config_data[1]~FF  (.D(1'b1), .CE(\uart_rx_inst/n1161 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx_inst/r_config_data [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(168)
    defparam \uart_rx_inst/r_config_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_config_data[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx_inst/r_config_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_config_data[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx_inst/r_config_data[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx_inst/r_config_data[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx_inst/r_config_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[1]~FF  (.D(rx_data[1]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \b[1]~FF .CLK_POLARITY = 1'b1;
    defparam \b[1]~FF .CE_POLARITY = 1'b1;
    defparam \b[1]~FF .SR_POLARITY = 1'b1;
    defparam \b[1]~FF .D_POLARITY = 1'b1;
    defparam \b[1]~FF .SR_SYNC = 1'b1;
    defparam \b[1]~FF .SR_VALUE = 1'b0;
    defparam \b[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[2]~FF  (.D(rx_data[2]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \b[2]~FF .CLK_POLARITY = 1'b1;
    defparam \b[2]~FF .CE_POLARITY = 1'b1;
    defparam \b[2]~FF .SR_POLARITY = 1'b1;
    defparam \b[2]~FF .D_POLARITY = 1'b1;
    defparam \b[2]~FF .SR_SYNC = 1'b1;
    defparam \b[2]~FF .SR_VALUE = 1'b0;
    defparam \b[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \b[3]~FF  (.D(rx_data[3]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(b[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \b[3]~FF .CLK_POLARITY = 1'b1;
    defparam \b[3]~FF .CE_POLARITY = 1'b1;
    defparam \b[3]~FF .SR_POLARITY = 1'b1;
    defparam \b[3]~FF .D_POLARITY = 1'b1;
    defparam \b[3]~FF .SR_SYNC = 1'b1;
    defparam \b[3]~FF .SR_VALUE = 1'b0;
    defparam \b[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \sum[1]~FF  (.D(n25[1]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(sum[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \sum[1]~FF .CLK_POLARITY = 1'b1;
    defparam \sum[1]~FF .CE_POLARITY = 1'b1;
    defparam \sum[1]~FF .SR_POLARITY = 1'b1;
    defparam \sum[1]~FF .D_POLARITY = 1'b1;
    defparam \sum[1]~FF .SR_SYNC = 1'b1;
    defparam \sum[1]~FF .SR_VALUE = 1'b0;
    defparam \sum[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \sum[2]~FF  (.D(n25[2]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(sum[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \sum[2]~FF .CLK_POLARITY = 1'b1;
    defparam \sum[2]~FF .CE_POLARITY = 1'b1;
    defparam \sum[2]~FF .SR_POLARITY = 1'b1;
    defparam \sum[2]~FF .D_POLARITY = 1'b1;
    defparam \sum[2]~FF .SR_SYNC = 1'b1;
    defparam \sum[2]~FF .SR_VALUE = 1'b0;
    defparam \sum[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \sum[3]~FF  (.D(n25[3]), .CE(add_flag), .CLK(\clk~O ), .SR(1'b0), 
           .Q(sum[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \sum[3]~FF .CLK_POLARITY = 1'b1;
    defparam \sum[3]~FF .CE_POLARITY = 1'b1;
    defparam \sum[3]~FF .SR_POLARITY = 1'b1;
    defparam \sum[3]~FF .D_POLARITY = 1'b1;
    defparam \sum[3]~FF .SR_SYNC = 1'b1;
    defparam \sum[3]~FF .SR_VALUE = 1'b0;
    defparam \sum[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[0]~FF  (.D(\uart_tx_inst/n1116 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_2~FF  (.D(\uart_tx_inst/n733 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(tx_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \tx_2~FF .CLK_POLARITY = 1'b1;
    defparam \tx_2~FF .CE_POLARITY = 1'b0;
    defparam \tx_2~FF .SR_POLARITY = 1'b1;
    defparam \tx_2~FF .D_POLARITY = 1'b0;
    defparam \tx_2~FF .SR_SYNC = 1'b1;
    defparam \tx_2~FF .SR_VALUE = 1'b0;
    defparam \tx_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[0]~FF  (.D(\uart_tx_inst/n1120 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[0]~FF  (.D(\uart_tx_inst/n1112 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_tx_inst/r_SM_Main [2]), .Q(\uart_tx_inst/r_SM_Main [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[1]~FF  (.D(\uart_tx_inst/n786 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[2]~FF  (.D(\uart_tx_inst/n789 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[3]~FF  (.D(\uart_tx_inst/n792 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[4]~FF  (.D(\uart_tx_inst/n795 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[5]~FF  (.D(\uart_tx_inst/n798 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[6]~FF  (.D(\uart_tx_inst/n801 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[7]~FF  (.D(\uart_tx_inst/n804 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[8]~FF  (.D(\uart_tx_inst/n807 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[9]~FF  (.D(\uart_tx_inst/n810 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[10]~FF  (.D(\uart_tx_inst/n813 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[11]~FF  (.D(\uart_tx_inst/n816 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[12]~FF  (.D(\uart_tx_inst/n819 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[13]~FF  (.D(\uart_tx_inst/n822 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[14]~FF  (.D(\uart_tx_inst/n825 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[15]~FF  (.D(\uart_tx_inst/n828 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[16]~FF  (.D(\uart_tx_inst/n831 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[17]~FF  (.D(\uart_tx_inst/n834 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[18]~FF  (.D(\uart_tx_inst/n837 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[19]~FF  (.D(\uart_tx_inst/n840 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[20]~FF  (.D(\uart_tx_inst/n843 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[21]~FF  (.D(\uart_tx_inst/n846 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[22]~FF  (.D(\uart_tx_inst/n849 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[23]~FF  (.D(\uart_tx_inst/n852 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[24]~FF  (.D(\uart_tx_inst/n855 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[25]~FF  (.D(\uart_tx_inst/n858 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[26]~FF  (.D(\uart_tx_inst/n861 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[27]~FF  (.D(\uart_tx_inst/n864 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[28]~FF  (.D(\uart_tx_inst/n867 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[29]~FF  (.D(\uart_tx_inst/n870 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[30]~FF  (.D(\uart_tx_inst/n873 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Clock_Count[31]~FF  (.D(\uart_tx_inst/n876 ), .CE(\uart_tx_inst/r_SM_Main [2]), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Clock_Count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Clock_Count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[1]~FF  (.D(\uart_tx_inst/n880 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Bit_Index[2]~FF  (.D(\uart_tx_inst/n884 ), .CE(ceg_net28), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Bit_Index [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_config_data[31]~FF  (.D(1'b1), .CE(\uart_tx_inst/n1032 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_config_data [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_config_data[31]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_config_data[31]~FF .CE_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_config_data[31]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_config_data[31]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_config_data[31]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_config_data[31]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_config_data[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[3]~FF  (.D(carry), .CE(\uart_tx_inst/n1224 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[4]~FF  (.D(sum[0]), .CE(\uart_tx_inst/n1224 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[5]~FF  (.D(sum[1]), .CE(\uart_tx_inst/n1224 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[6]~FF  (.D(sum[2]), .CE(\uart_tx_inst/n1224 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_Tx_Data[7]~FF  (.D(sum[3]), .CE(\uart_tx_inst/n1224 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx_inst/r_Tx_Data [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_Tx_Data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[1]~FF  (.D(\uart_tx_inst/n779 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_tx_inst/r_SM_Main [2]), .Q(\uart_tx_inst/r_SM_Main [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx_inst/r_SM_Main[2]~FF  (.D(\uart_tx_inst/n50 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\uart_tx_inst/n1206 ), .Q(\uart_tx_inst/r_SM_Main [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam \uart_tx_inst/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx_inst/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[1]~FF  (.D(rx_data[5]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \a[1]~FF .CLK_POLARITY = 1'b1;
    defparam \a[1]~FF .CE_POLARITY = 1'b1;
    defparam \a[1]~FF .SR_POLARITY = 1'b1;
    defparam \a[1]~FF .D_POLARITY = 1'b1;
    defparam \a[1]~FF .SR_SYNC = 1'b1;
    defparam \a[1]~FF .SR_VALUE = 1'b0;
    defparam \a[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[2]~FF  (.D(rx_data[6]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \a[2]~FF .CLK_POLARITY = 1'b1;
    defparam \a[2]~FF .CE_POLARITY = 1'b1;
    defparam \a[2]~FF .SR_POLARITY = 1'b1;
    defparam \a[2]~FF .D_POLARITY = 1'b1;
    defparam \a[2]~FF .SR_SYNC = 1'b1;
    defparam \a[2]~FF .SR_VALUE = 1'b0;
    defparam \a[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \a[3]~FF  (.D(rx_data[7]), .CE(rx_ready), .CLK(\clk~O ), .SR(1'b0), 
           .Q(a[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(38)
    defparam \a[3]~FF .CLK_POLARITY = 1'b1;
    defparam \a[3]~FF .CE_POLARITY = 1'b1;
    defparam \a[3]~FF .SR_POLARITY = 1'b1;
    defparam \a[3]~FF .D_POLARITY = 1'b1;
    defparam \a[3]~FF .SR_SYNC = 1'b1;
    defparam \a[3]~FF .SR_VALUE = 1'b0;
    defparam \a[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n999 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1000 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1001 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/skip_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1757 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3659)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [0]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3688)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n1975 [0]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [0]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2194 [0]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state [0]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3770)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/n2545 ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4080)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n2558 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n2545 ), .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4080)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(rx_ready), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n2558 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(rx_data[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3447 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3447 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr [0]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr [64]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1055 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3621)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[8]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[9]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[10]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[11]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[12]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[13]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[14]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[15]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[16]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[17]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[18]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[19]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[20]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[21]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[22]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[23]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[24]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[25]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[26]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[27]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[28]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[29]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[30]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[31]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[32]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[33]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[34]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[35]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[36]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[37]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[38]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[39]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[40]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[41]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[42]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[43]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[44]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[45]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[46]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[47]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[48]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[49]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[50]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[51]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[52]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[53]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[54]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[55]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[56]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[57]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[58]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[59]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[60]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[61]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[62]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/skip_count[63]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1572 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/skip_count [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3631)
    defparam \edb_top_inst/la0/skip_count[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/skip_count[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/la0/n1705 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3644)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [1]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [2]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [3]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [4]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [5]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [6]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [7]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [8]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [9]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [10]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [11]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [12]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [13]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [14]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [15]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [16]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [17]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [18]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [19]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [20]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [21]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [22]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [23]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter [24]), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3678)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3688)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3688)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3688)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n1975 [1]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n1975 [2]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n1975 [3]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n1975 [4]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n1975 [5]), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [1]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [2]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [3]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [4]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [5]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [6]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [7]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [8]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [9]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [10]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [11]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [12]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [13]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [14]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter [15]), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3715)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2194 [1]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2194 [2]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2194 [3]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2194 [4]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2194 [5]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2194 [6]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2194 [7]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2194 [8]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2194 [9]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2194 [10]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2194 [11]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2194 [12]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2194 [13]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2194 [14]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2194 [15]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2194 [16]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2194 [17]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2194 [18]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2194 [19]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2194 [20]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2194 [21]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2194 [22]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2194 [23]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2194 [24]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2194 [25]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2194 [26]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2194 [27]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2194 [28]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2194 [29]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2194 [30]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2194 [31]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2194 [32]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2194 [33]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2194 [34]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2194 [35]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2194 [36]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2194 [37]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2194 [38]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2194 [39]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2194 [40]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2194 [41]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2194 [42]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2194 [43]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2194 [44]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2194 [45]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2194 [46]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2194 [47]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2194 [48]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2194 [49]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2194 [50]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2194 [51]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2194 [52]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2194 [53]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2194 [54]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2194 [55]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2194 [56]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2194 [57]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2194 [58]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2194 [59]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2194 [60]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2194 [61]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2194 [62]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2194 [63]), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3728)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state [1]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3770)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state [2]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3770)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state [3]), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3770)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [0]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [1]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [2]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [3]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [4]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [5]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [6]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [7]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [8]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [9]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [10]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [11]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [12]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [13]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [14]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [15]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [16]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [17]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [18]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [19]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [20]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [21]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [22]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [23]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [24]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [25]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [26]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [27]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [28]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [29]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [30]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n118 [31]), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(240)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n2558 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF  (.D(rx_data[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF  (.D(rx_data[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF  (.D(rx_data[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF  (.D(rx_data[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF  (.D(rx_data[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF  (.D(rx_data[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF  (.D(rx_data[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4107)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5516)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5577)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5516)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3447 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n3462 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/la0/n3660 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5628)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n29 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5758)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[8]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1 [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4404)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4416)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [0]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/ts_trigger~FF  (.D(1'b1), .CE(\edb_top_inst/la0/trigger_skipper_n/n468 ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), .Q(\edb_top_inst/la0/ts_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/ts_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/ts_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [1]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [2]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [3]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [4]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [5]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [6]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [7]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [8]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [9]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [10]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [11]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [12]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [13]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [14]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [15]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [16]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [17]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [18]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [19]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [20]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [21]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [22]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [23]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [24]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [25]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [26]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [27]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [28]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [29]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [30]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [31]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [32]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [33]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [34]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [35]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [36]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [37]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [38]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [39]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [40]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [41]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [42]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [43]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [44]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [45]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [46]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [47]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [48]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [49]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [50]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [51]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [52]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [53]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [54]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [55]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [56]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [57]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [58]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [59]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [60]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [61]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [62]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF  (.D(\edb_top_inst/la0/trigger_skipper_n/n138 [63]), 
           .CE(\edb_top_inst/la0/tu_trigger ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/ts_resetn ), 
           .Q(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5833)
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5244)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5044)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5044)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5044)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/ts_resetn~FF  (.D(\edb_top_inst/la0/la_biu_inst/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/ts_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5044)
    defparam \edb_top_inst/la0/ts_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/ts_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5265)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5280)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5280)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5280)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5290)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5303)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5303)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5303)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1249 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/n1832 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5427)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1214 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n5970 ), .Q(\edb_top_inst/la0/la_biu_inst/curr_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5244)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5244)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5244)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5044)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n335 ), 
           .CE(\edb_top_inst/ceg_net18 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5315)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter [15]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter [16]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter [17]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter [18]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter [19]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter [20]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter [21]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter [22]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter [23]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter [24]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n335 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5325)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1248 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5334)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state [1]), 
           .CE(\edb_top_inst/ceg_net24 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5427)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt [0]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1839 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1839 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [1]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [2]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [3]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [4]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [5]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [6]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [7]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [8]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [9]), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 [1]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [2]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [3]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [4]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [5]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [6]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [7]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [8]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [9]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [10]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4736)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4558)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n110 [1]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [2]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [3]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [4]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [5]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [6]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [7]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [8]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [9]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [10]), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4653)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr [65]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr [66]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr [67]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr [68]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr [69]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr [70]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr [71]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr [72]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr [73]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr [74]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr [75]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr [76]), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3561)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/la0/n971 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3611)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(311)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr [1]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(311)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(311)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(311)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr [2]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr [3]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr [4]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr [5]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr [6]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr [7]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr [8]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr [9]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr [10]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr [11]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr [12]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr [13]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr [14]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr [15]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr [16]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr [17]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr [18]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr [19]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr [20]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr [21]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr [22]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr [23]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr [24]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr [25]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr [26]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr [27]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr [28]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr [29]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr [30]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr [31]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr [32]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr [33]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr [34]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr [35]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr [36]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr [37]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr [38]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr [39]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr [40]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr [41]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr [42]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr [43]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr [44]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr [45]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr [46]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr [47]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr [48]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr [49]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr [50]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr [51]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr [52]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr [53]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr [54]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr [55]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr [56]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr [57]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr [58]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr [59]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr [60]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr [61]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr [62]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr [63]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr [64]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr [65]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr [66]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr [67]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr [68]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr [69]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr [70]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr [71]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr [72]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr [73]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr [74]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr [75]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr [76]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr [77]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr [78]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr [79]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr [80]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr [81]), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr [81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(304)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \edb_top_inst/LUT__2994  (.I0(\edb_top_inst/la0/crc_data_out [29]), 
            .I1(\edb_top_inst/edb_user_dr [79]), .I2(\edb_top_inst/la0/crc_data_out [30]), 
            .I3(\edb_top_inst/edb_user_dr [80]), .O(\edb_top_inst/n1407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2994 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2995  (.I0(\edb_top_inst/la0/crc_data_out [27]), 
            .I1(\edb_top_inst/edb_user_dr [77]), .I2(\edb_top_inst/la0/crc_data_out [28]), 
            .I3(\edb_top_inst/edb_user_dr [78]), .O(\edb_top_inst/n1408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2995 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2996  (.I0(\edb_top_inst/la0/crc_data_out [25]), 
            .I1(\edb_top_inst/edb_user_dr [75]), .I2(\edb_top_inst/la0/crc_data_out [26]), 
            .I3(\edb_top_inst/edb_user_dr [76]), .O(\edb_top_inst/n1409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2996 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2997  (.I0(\edb_top_inst/n1406 ), .I1(\edb_top_inst/n1407 ), 
            .I2(\edb_top_inst/n1408 ), .I3(\edb_top_inst/n1409 ), .O(\edb_top_inst/n1410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2997 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2998  (.I0(\edb_top_inst/la0/crc_data_out [21]), 
            .I1(\edb_top_inst/edb_user_dr [71]), .I2(\edb_top_inst/la0/crc_data_out [22]), 
            .I3(\edb_top_inst/edb_user_dr [72]), .O(\edb_top_inst/n1411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2998 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2999  (.I0(\edb_top_inst/la0/crc_data_out [16]), 
            .I1(\edb_top_inst/edb_user_dr [66]), .I2(\edb_top_inst/la0/crc_data_out [23]), 
            .I3(\edb_top_inst/edb_user_dr [73]), .O(\edb_top_inst/n1412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2999 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3000  (.I0(\edb_top_inst/la0/crc_data_out [19]), 
            .I1(\edb_top_inst/edb_user_dr [69]), .I2(\edb_top_inst/la0/crc_data_out [20]), 
            .I3(\edb_top_inst/edb_user_dr [70]), .O(\edb_top_inst/n1413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3000 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3001  (.I0(\edb_top_inst/la0/crc_data_out [17]), 
            .I1(\edb_top_inst/edb_user_dr [67]), .I2(\edb_top_inst/la0/crc_data_out [18]), 
            .I3(\edb_top_inst/edb_user_dr [68]), .O(\edb_top_inst/n1414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3001 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3002  (.I0(\edb_top_inst/n1411 ), .I1(\edb_top_inst/n1412 ), 
            .I2(\edb_top_inst/n1413 ), .I3(\edb_top_inst/n1414 ), .O(\edb_top_inst/n1415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3002 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3003  (.I0(\edb_top_inst/la0/crc_data_out [8]), 
            .I1(\edb_top_inst/edb_user_dr [58]), .I2(\edb_top_inst/la0/crc_data_out [9]), 
            .I3(\edb_top_inst/edb_user_dr [59]), .O(\edb_top_inst/n1416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3003 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3004  (.I0(\edb_top_inst/la0/crc_data_out [10]), 
            .I1(\edb_top_inst/edb_user_dr [60]), .I2(\edb_top_inst/la0/crc_data_out [11]), 
            .I3(\edb_top_inst/edb_user_dr [61]), .O(\edb_top_inst/n1417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3004 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3005  (.I0(\edb_top_inst/la0/crc_data_out [12]), 
            .I1(\edb_top_inst/edb_user_dr [62]), .I2(\edb_top_inst/la0/crc_data_out [13]), 
            .I3(\edb_top_inst/edb_user_dr [63]), .O(\edb_top_inst/n1418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3005 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3006  (.I0(\edb_top_inst/la0/crc_data_out [7]), 
            .I1(\edb_top_inst/edb_user_dr [57]), .I2(\edb_top_inst/la0/crc_data_out [14]), 
            .I3(\edb_top_inst/edb_user_dr [64]), .O(\edb_top_inst/n1419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3006 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3007  (.I0(\edb_top_inst/n1416 ), .I1(\edb_top_inst/n1417 ), 
            .I2(\edb_top_inst/n1418 ), .I3(\edb_top_inst/n1419 ), .O(\edb_top_inst/n1420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3007 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3008  (.I0(\edb_top_inst/la0/crc_data_out [0]), 
            .I1(\edb_top_inst/edb_user_dr [50]), .I2(\edb_top_inst/la0/crc_data_out [1]), 
            .I3(\edb_top_inst/edb_user_dr [51]), .O(\edb_top_inst/n1421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3008 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3009  (.I0(\edb_top_inst/la0/crc_data_out [2]), 
            .I1(\edb_top_inst/edb_user_dr [52]), .I2(\edb_top_inst/la0/crc_data_out [3]), 
            .I3(\edb_top_inst/edb_user_dr [53]), .O(\edb_top_inst/n1422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3009 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3010  (.I0(\edb_top_inst/la0/crc_data_out [6]), 
            .I1(\edb_top_inst/edb_user_dr [56]), .I2(\edb_top_inst/la0/crc_data_out [15]), 
            .I3(\edb_top_inst/edb_user_dr [65]), .O(\edb_top_inst/n1423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3010 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3011  (.I0(\edb_top_inst/la0/crc_data_out [4]), 
            .I1(\edb_top_inst/edb_user_dr [54]), .I2(\edb_top_inst/la0/crc_data_out [5]), 
            .I3(\edb_top_inst/edb_user_dr [55]), .O(\edb_top_inst/n1424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3011 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3012  (.I0(\edb_top_inst/n1421 ), .I1(\edb_top_inst/n1422 ), 
            .I2(\edb_top_inst/n1423 ), .I3(\edb_top_inst/n1424 ), .O(\edb_top_inst/n1425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3012 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3013  (.I0(\edb_top_inst/n1410 ), .I1(\edb_top_inst/n1415 ), 
            .I2(\edb_top_inst/n1420 ), .I3(\edb_top_inst/n1425 ), .O(\edb_top_inst/n1426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3013 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3014  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/crc_data_out [0]), .I2(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n1427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3014 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3015  (.I0(\edb_top_inst/n1427 ), .I1(\edb_top_inst/n1426 ), 
            .I2(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n1428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3015 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3016  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n1429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3016 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3017  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n1430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3017 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3018  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg [0]), .I2(\edb_top_inst/n1429 ), 
            .I3(\edb_top_inst/n1430 ), .O(\edb_top_inst/n1431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3018 .LUTMASK = 16'h5333;
    EFX_LUT4 \edb_top_inst/LUT__3019  (.I0(\edb_top_inst/la0/bit_count [3]), 
            .I1(\edb_top_inst/la0/bit_count [4]), .I2(\edb_top_inst/la0/bit_count [5]), 
            .O(\edb_top_inst/n1432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3019 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3020  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/la0/bit_count [1]), .I2(\edb_top_inst/la0/bit_count [2]), 
            .O(\edb_top_inst/n1433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3020 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3021  (.I0(\edb_top_inst/la0/word_count [8]), 
            .I1(\edb_top_inst/la0/word_count [9]), .I2(\edb_top_inst/la0/word_count [10]), 
            .I3(\edb_top_inst/la0/word_count [11]), .O(\edb_top_inst/n1434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3021 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3022  (.I0(\edb_top_inst/la0/word_count [4]), 
            .I1(\edb_top_inst/la0/word_count [5]), .I2(\edb_top_inst/la0/word_count [6]), 
            .I3(\edb_top_inst/la0/word_count [7]), .O(\edb_top_inst/n1435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3022 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3023  (.I0(\edb_top_inst/la0/word_count [0]), 
            .I1(\edb_top_inst/la0/word_count [1]), .I2(\edb_top_inst/la0/word_count [2]), 
            .I3(\edb_top_inst/la0/word_count [3]), .O(\edb_top_inst/n1436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3023 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3024  (.I0(\edb_top_inst/la0/word_count [12]), 
            .I1(\edb_top_inst/la0/word_count [13]), .I2(\edb_top_inst/la0/word_count [14]), 
            .I3(\edb_top_inst/la0/word_count [15]), .O(\edb_top_inst/n1437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3024 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3025  (.I0(\edb_top_inst/n1434 ), .I1(\edb_top_inst/n1435 ), 
            .I2(\edb_top_inst/n1436 ), .I3(\edb_top_inst/n1437 ), .O(\edb_top_inst/n1438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3025 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3026  (.I0(\edb_top_inst/n1433 ), .I1(\edb_top_inst/n1432 ), 
            .I2(\edb_top_inst/n1438 ), .I3(\edb_top_inst/la0/module_state [1]), 
            .O(\edb_top_inst/n1439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3026 .LUTMASK = 16'h77f0;
    EFX_LUT4 \edb_top_inst/LUT__3027  (.I0(\edb_top_inst/n1439 ), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(jtag_inst1_UPDATE), .O(\edb_top_inst/n1440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3027 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__3028  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg [1]), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg [2]), .I2(\edb_top_inst/debug_hub_inst/module_id_reg [3]), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg [0]), .O(\edb_top_inst/n1441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3028 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3029  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n1442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3029 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3030  (.I0(\edb_top_inst/n1441 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n1442 ), .I3(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n1443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3030 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__3031  (.I0(\edb_top_inst/edb_user_dr [77]), 
            .I1(\edb_top_inst/edb_user_dr [78]), .I2(\edb_top_inst/edb_user_dr [79]), 
            .I3(\edb_top_inst/edb_user_dr [80]), .O(\edb_top_inst/n1444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3031 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__3032  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n1445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3032 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3033  (.I0(\edb_top_inst/edb_user_dr [81]), 
            .I1(jtag_inst1_UPDATE), .O(\edb_top_inst/n1446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3033 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3034  (.I0(\edb_top_inst/n1444 ), .I1(\edb_top_inst/n1445 ), 
            .I2(\edb_top_inst/n1441 ), .I3(\edb_top_inst/n1446 ), .O(\edb_top_inst/n1447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3034 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3035  (.I0(\edb_top_inst/n1443 ), .I1(\edb_top_inst/la0/module_state [1]), 
            .I2(\edb_top_inst/n1447 ), .O(\edb_top_inst/n1448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3035 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3036  (.I0(\edb_top_inst/n1448 ), .I1(\edb_top_inst/n1440 ), 
            .I2(\edb_top_inst/la0/module_state [2]), .I3(\edb_top_inst/la0/module_state [3]), 
            .O(\edb_top_inst/n1449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3036 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__3037  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n1450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3037 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3038  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/n1449 ), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/n1450 ), .O(\edb_top_inst/n1451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3038 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__3039  (.I0(\edb_top_inst/n1431 ), .I1(\edb_top_inst/n1428 ), 
            .I2(\edb_top_inst/n1451 ), .I3(\edb_top_inst/n1441 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3039 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3040  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [40]), .O(\edb_top_inst/la0/n999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3040 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3041  (.I0(\edb_top_inst/edb_user_dr [66]), 
            .I1(\edb_top_inst/edb_user_dr [67]), .I2(\edb_top_inst/edb_user_dr [68]), 
            .I3(\edb_top_inst/edb_user_dr [69]), .O(\edb_top_inst/n1452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3041 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3042  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n1452 ), 
            .O(\edb_top_inst/n1453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3042 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3043  (.I0(\edb_top_inst/edb_user_dr [74]), 
            .I1(\edb_top_inst/edb_user_dr [75]), .I2(\edb_top_inst/edb_user_dr [76]), 
            .I3(\edb_top_inst/edb_user_dr [79]), .O(\edb_top_inst/n1454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3043 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3044  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .I2(\edb_top_inst/la0/module_state [2]), 
            .I3(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n1455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3044 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3045  (.I0(\edb_top_inst/edb_user_dr [78]), 
            .I1(\edb_top_inst/edb_user_dr [77]), .I2(\edb_top_inst/edb_user_dr [80]), 
            .O(\edb_top_inst/n1456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3045 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3046  (.I0(\edb_top_inst/n1441 ), .I1(\edb_top_inst/n1446 ), 
            .I2(\edb_top_inst/n1455 ), .I3(\edb_top_inst/n1456 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3046 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3047  (.I0(\edb_top_inst/edb_user_dr [70]), 
            .I1(\edb_top_inst/edb_user_dr [73]), .I2(\edb_top_inst/n1454 ), 
            .I3(\edb_top_inst/la0/regsel_ld_en ), .O(\edb_top_inst/n1457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3047 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3048  (.I0(\edb_top_inst/edb_user_dr [72]), 
            .I1(\edb_top_inst/n1457 ), .O(\edb_top_inst/n1458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3048 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3049  (.I0(\edb_top_inst/edb_user_dr [71]), 
            .I1(\edb_top_inst/n1458 ), .O(\edb_top_inst/n1459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3049 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3050  (.I0(\edb_top_inst/n1453 ), .I1(\edb_top_inst/n1459 ), 
            .O(\edb_top_inst/la0/n971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3050 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3051  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/la0/n971 ), .O(\edb_top_inst/ceg_net2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3051 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3052  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [41]), .O(\edb_top_inst/la0/n1000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3052 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3053  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr [42]), .O(\edb_top_inst/la0/n1001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3053 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3054  (.I0(\edb_top_inst/edb_user_dr [65]), 
            .I1(\edb_top_inst/edb_user_dr [64]), .I2(\edb_top_inst/n1452 ), 
            .I3(\edb_top_inst/n1459 ), .O(\edb_top_inst/la0/n1055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3054 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3055  (.I0(\edb_top_inst/edb_user_dr [66]), 
            .I1(\edb_top_inst/edb_user_dr [68]), .I2(\edb_top_inst/edb_user_dr [69]), 
            .I3(\edb_top_inst/edb_user_dr [67]), .O(\edb_top_inst/n1460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3055 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3056  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n1459 ), 
            .I3(\edb_top_inst/n1460 ), .O(\edb_top_inst/la0/n1572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3056 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3057  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n1452 ), 
            .I3(\edb_top_inst/n1459 ), .O(\edb_top_inst/la0/n1705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3057 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3058  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/edb_user_dr [68]), 
            .I3(\edb_top_inst/edb_user_dr [69]), .O(\edb_top_inst/n1461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3058 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3059  (.I0(\edb_top_inst/edb_user_dr [67]), 
            .I1(\edb_top_inst/edb_user_dr [66]), .I2(\edb_top_inst/edb_user_dr [63]), 
            .I3(\edb_top_inst/n1461 ), .O(\edb_top_inst/n1462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3059 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3060  (.I0(\edb_top_inst/n1459 ), .I1(\edb_top_inst/n1462 ), 
            .O(\edb_top_inst/la0/n1757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3060 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3061  (.I0(\edb_top_inst/la0/address_counter [4]), 
            .I1(\edb_top_inst/la0/address_counter [5]), .I2(\edb_top_inst/la0/address_counter [6]), 
            .I3(\edb_top_inst/la0/address_counter [7]), .O(\edb_top_inst/n1463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3061 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3062  (.I0(\edb_top_inst/la0/address_counter [0]), 
            .I1(\edb_top_inst/la0/address_counter [1]), .I2(\edb_top_inst/la0/address_counter [2]), 
            .I3(\edb_top_inst/la0/address_counter [3]), .O(\edb_top_inst/n1464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3062 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3063  (.I0(\edb_top_inst/la0/address_counter [8]), 
            .I1(\edb_top_inst/la0/address_counter [9]), .I2(\edb_top_inst/la0/address_counter [10]), 
            .I3(\edb_top_inst/la0/address_counter [11]), .O(\edb_top_inst/n1465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3063 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3064  (.I0(\edb_top_inst/la0/address_counter [12]), 
            .I1(\edb_top_inst/la0/address_counter [13]), .I2(\edb_top_inst/la0/address_counter [14]), 
            .O(\edb_top_inst/n1466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3064 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3065  (.I0(\edb_top_inst/n1463 ), .I1(\edb_top_inst/n1464 ), 
            .I2(\edb_top_inst/n1465 ), .I3(\edb_top_inst/n1466 ), .O(\edb_top_inst/n1467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3065 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3066  (.I0(\edb_top_inst/n1467 ), .I1(\edb_top_inst/la0/n1814 [0]), 
            .I2(\edb_top_inst/edb_user_dr [45]), .I3(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3066 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3067  (.I0(\edb_top_inst/n1447 ), .I1(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3067 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3068  (.I0(\edb_top_inst/n1445 ), .I1(\edb_top_inst/la0/module_state [3]), 
            .I2(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n1468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3068 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3069  (.I0(\edb_top_inst/la0/word_count [1]), 
            .I1(\edb_top_inst/la0/word_count [2]), .I2(\edb_top_inst/la0/word_count [3]), 
            .O(\edb_top_inst/n1469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3069 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3070  (.I0(\edb_top_inst/n1434 ), .I1(\edb_top_inst/n1435 ), 
            .I2(\edb_top_inst/n1437 ), .I3(\edb_top_inst/n1469 ), .O(\edb_top_inst/n1470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3070 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3071  (.I0(\edb_top_inst/la0/opcode [3]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [0]), .O(\edb_top_inst/la0/n595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3071 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3072  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [3]), .O(\edb_top_inst/la0/n596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3072 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3073  (.I0(\edb_top_inst/la0/n595 ), .I1(\edb_top_inst/la0/bit_count [5]), 
            .I2(\edb_top_inst/la0/n596 ), .I3(\edb_top_inst/la0/bit_count [4]), 
            .O(\edb_top_inst/n1471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3073 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__3074  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [1]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [3]), .O(\edb_top_inst/n1472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3074 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__3075  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/la0/bit_count [1]), .I2(\edb_top_inst/la0/bit_count [2]), 
            .I3(\edb_top_inst/n1472 ), .O(\edb_top_inst/n1473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3075 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__3076  (.I0(\edb_top_inst/la0/opcode [1]), 
            .I1(\edb_top_inst/la0/opcode [3]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [0]), .O(\edb_top_inst/la0/n593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3076 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3077  (.I0(\edb_top_inst/n1472 ), .I1(\edb_top_inst/la0/n593 ), 
            .I2(\edb_top_inst/la0/bit_count [3]), .O(\edb_top_inst/n1474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3077 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__3078  (.I0(\edb_top_inst/n1471 ), .I1(\edb_top_inst/n1473 ), 
            .I2(\edb_top_inst/n1474 ), .O(\edb_top_inst/n1475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3078 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3079  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/la0/module_state [1]), .I2(\edb_top_inst/n1475 ), 
            .O(\edb_top_inst/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3079 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__3080  (.I0(\edb_top_inst/n1470 ), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(\edb_top_inst/la0/module_state [3]), .I3(\edb_top_inst/n1476 ), 
            .O(\edb_top_inst/n1477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3080 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__3081  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/n1438 ), .I2(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n1478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3081 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3082  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/n1429 ), .I3(\edb_top_inst/n1430 ), .O(\edb_top_inst/n1479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3082 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3083  (.I0(\edb_top_inst/n1479 ), .I1(\edb_top_inst/n1470 ), 
            .I2(\edb_top_inst/n1430 ), .O(\edb_top_inst/n1480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3083 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__3084  (.I0(\edb_top_inst/n1478 ), .I1(\edb_top_inst/n1480 ), 
            .I2(\edb_top_inst/n1468 ), .I3(\edb_top_inst/n1477 ), .O(\edb_top_inst/n1481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3084 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__3085  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n1481 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3085 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3086  (.I0(\edb_top_inst/n1447 ), .I1(\edb_top_inst/la0/module_state [3]), 
            .I2(\edb_top_inst/n1445 ), .O(\edb_top_inst/n1482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3086 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__3087  (.I0(\edb_top_inst/la0/module_state [2]), 
            .I1(\edb_top_inst/n1479 ), .I2(\edb_top_inst/n1482 ), .O(\edb_top_inst/n1483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3087 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3088  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/n1476 ), .I2(\edb_top_inst/la0/module_state [2]), 
            .I3(\edb_top_inst/n1483 ), .O(\edb_top_inst/n1484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3088 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__3089  (.I0(\edb_top_inst/la0/bit_count [0]), 
            .I1(\edb_top_inst/n1484 ), .O(\edb_top_inst/la0/n1975 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3089 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3090  (.I0(\edb_top_inst/n1438 ), .I1(\edb_top_inst/n1475 ), 
            .O(\edb_top_inst/n1485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3090 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3091  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/n1485 ), 
            .O(\edb_top_inst/n1486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3091 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__3092  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/edb_user_dr [81]), 
            .O(\edb_top_inst/n1487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3092 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3093  (.I0(\edb_top_inst/n1487 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n1478 ), .I3(\edb_top_inst/n1441 ), .O(\edb_top_inst/n1488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbaf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3093 .LUTMASK = 16'hbaf0;
    EFX_LUT4 \edb_top_inst/LUT__3094  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n1489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3094 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3095  (.I0(\edb_top_inst/n1488 ), .I1(\edb_top_inst/n1486 ), 
            .I2(\edb_top_inst/n1489 ), .I3(\edb_top_inst/n1449 ), .O(\edb_top_inst/la0/module_next_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3095 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__3096  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/n1489 ), .O(\edb_top_inst/n1490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3096 .LUTMASK = 16'he300;
    EFX_LUT4 \edb_top_inst/LUT__3097  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/module_state [0]), 
            .I2(\edb_top_inst/n1490 ), .I3(\edb_top_inst/n1450 ), .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3097 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__3098  (.I0(\edb_top_inst/edb_user_dr [29]), 
            .I1(\edb_top_inst/la0/word_count [0]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_word_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3098 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__3099  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/n1475 ), .I2(\edb_top_inst/la0/module_state [0]), 
            .I3(\edb_top_inst/la0/module_state [1]), .O(\edb_top_inst/n1491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3099 .LUTMASK = 16'h35f3;
    EFX_LUT4 \edb_top_inst/LUT__3100  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/n1491 ), .I2(\edb_top_inst/la0/module_state [2]), 
            .I3(\edb_top_inst/n1483 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3100 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__3101  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/n1492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3101 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__3102  (.I0(\edb_top_inst/la0/internal_register_select [9]), 
            .I1(\edb_top_inst/la0/internal_register_select [10]), .I2(\edb_top_inst/la0/internal_register_select [11]), 
            .I3(\edb_top_inst/la0/internal_register_select [12]), .O(\edb_top_inst/n1493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3102 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3103  (.I0(\edb_top_inst/la0/internal_register_select [2]), 
            .I1(\edb_top_inst/la0/internal_register_select [6]), .I2(\edb_top_inst/la0/internal_register_select [7]), 
            .I3(\edb_top_inst/la0/internal_register_select [8]), .O(\edb_top_inst/n1494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3103 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3104  (.I0(\edb_top_inst/n1493 ), .I1(\edb_top_inst/n1494 ), 
            .O(\edb_top_inst/n1495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3104 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3105  (.I0(\edb_top_inst/la0/internal_register_select [4]), 
            .I1(\edb_top_inst/la0/internal_register_select [5]), .O(\edb_top_inst/n1496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3105 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3106  (.I0(\edb_top_inst/la0/internal_register_select [1]), 
            .I1(\edb_top_inst/n1495 ), .I2(\edb_top_inst/n1496 ), .O(\edb_top_inst/n1497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3106 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3107  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/n1497 ), .O(\edb_top_inst/n1498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3107 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3108  (.I0(\edb_top_inst/n1492 ), .I1(\edb_top_inst/la0/la_trig_mask [0]), 
            .I2(\edb_top_inst/la0/internal_register_select [0]), .I3(\edb_top_inst/n1498 ), 
            .O(\edb_top_inst/n1499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3108 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3109  (.I0(\edb_top_inst/la0/internal_register_select [3]), 
            .I1(\edb_top_inst/n1496 ), .O(\edb_top_inst/n1500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3109 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3110  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/la0/internal_register_select [1]), .I2(\edb_top_inst/n1495 ), 
            .I3(\edb_top_inst/n1500 ), .O(\edb_top_inst/n1501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3110 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3111  (.I0(\edb_top_inst/la0/internal_register_select [1]), 
            .I1(\edb_top_inst/la0/internal_register_select [3]), .I2(\edb_top_inst/n1495 ), 
            .I3(\edb_top_inst/n1496 ), .O(\edb_top_inst/n1502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3111 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3112  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3112 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3113  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [0]), 
            .I2(\edb_top_inst/n1503 ), .O(\edb_top_inst/n1504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3113 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3114  (.I0(\edb_top_inst/n1489 ), .I1(\edb_top_inst/n1475 ), 
            .I2(\edb_top_inst/n1445 ), .I3(\edb_top_inst/n1479 ), .O(\edb_top_inst/n1505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3114 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__3115  (.I0(\edb_top_inst/n1499 ), .I1(\edb_top_inst/n1504 ), 
            .I2(\edb_top_inst/la0/data_from_biu [0]), .I3(\edb_top_inst/n1505 ), 
            .O(\edb_top_inst/n1506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3115 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3116  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n1441 ), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/n1507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3116 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3117  (.I0(\edb_top_inst/n1507 ), .I1(\edb_top_inst/n1505 ), 
            .O(\edb_top_inst/n1508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3117 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3118  (.I0(\edb_top_inst/n1506 ), .I1(\edb_top_inst/la0/data_out_shift_reg [1]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3118 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3119  (.I0(\edb_top_inst/n1441 ), .I1(jtag_inst1_SHIFT), 
            .I2(\edb_top_inst/la0/module_state [2]), .O(\edb_top_inst/n1509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3119 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3120  (.I0(\edb_top_inst/la0/module_state [3]), 
            .I1(\edb_top_inst/n1509 ), .I2(\edb_top_inst/n1445 ), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/ceg_net8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3120 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__3121  (.I0(jtag_inst1_RESET), .I1(\edb_top_inst/la0/la_soft_reset_in ), 
            .O(\edb_top_inst/la0/n2545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3121 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3122  (.I0(\edb_top_inst/edb_user_dr [71]), 
            .I1(\edb_top_inst/n1453 ), .I2(\edb_top_inst/n1458 ), .O(\edb_top_inst/la0/n2558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3122 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3123  (.I0(\edb_top_inst/edb_user_dr [71]), 
            .I1(\edb_top_inst/edb_user_dr [72]), .I2(\edb_top_inst/n1457 ), 
            .O(\edb_top_inst/n1510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3123 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3124  (.I0(\edb_top_inst/n1453 ), .I1(\edb_top_inst/n1510 ), 
            .O(\edb_top_inst/la0/n3447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3124 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3125  (.I0(\edb_top_inst/edb_user_dr [65]), 
            .I1(\edb_top_inst/edb_user_dr [64]), .I2(\edb_top_inst/n1452 ), 
            .I3(\edb_top_inst/n1510 ), .O(\edb_top_inst/la0/n3462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3125 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3126  (.I0(\edb_top_inst/edb_user_dr [64]), 
            .I1(\edb_top_inst/edb_user_dr [65]), .I2(\edb_top_inst/n1452 ), 
            .I3(\edb_top_inst/n1510 ), .O(\edb_top_inst/la0/n3660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3126 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3127  (.I0(\edb_top_inst/n1467 ), .I1(\edb_top_inst/la0/n1814 [1]), 
            .I2(\edb_top_inst/edb_user_dr [46]), .I3(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3127 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3128  (.I0(\edb_top_inst/n1467 ), .I1(\edb_top_inst/la0/n1814 [2]), 
            .I2(\edb_top_inst/edb_user_dr [47]), .I3(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3128 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3129  (.I0(\edb_top_inst/n1467 ), .I1(\edb_top_inst/la0/n1814 [3]), 
            .I2(\edb_top_inst/edb_user_dr [48]), .I3(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3129 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3130  (.I0(\edb_top_inst/edb_user_dr [49]), 
            .I1(\edb_top_inst/la0/n1814 [4]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3130 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3131  (.I0(\edb_top_inst/edb_user_dr [50]), 
            .I1(\edb_top_inst/la0/n1814 [5]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3131 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3132  (.I0(\edb_top_inst/edb_user_dr [51]), 
            .I1(\edb_top_inst/la0/n1814 [6]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3132 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3133  (.I0(\edb_top_inst/edb_user_dr [52]), 
            .I1(\edb_top_inst/la0/n1814 [7]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3133 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3134  (.I0(\edb_top_inst/edb_user_dr [53]), 
            .I1(\edb_top_inst/la0/n1814 [8]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3134 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3135  (.I0(\edb_top_inst/edb_user_dr [54]), 
            .I1(\edb_top_inst/la0/n1814 [9]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3135 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3136  (.I0(\edb_top_inst/edb_user_dr [55]), 
            .I1(\edb_top_inst/la0/n1814 [10]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3136 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3137  (.I0(\edb_top_inst/edb_user_dr [56]), 
            .I1(\edb_top_inst/la0/n1814 [11]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3137 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3138  (.I0(\edb_top_inst/edb_user_dr [57]), 
            .I1(\edb_top_inst/la0/n1814 [12]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3138 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3139  (.I0(\edb_top_inst/edb_user_dr [58]), 
            .I1(\edb_top_inst/la0/n1814 [13]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3139 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3140  (.I0(\edb_top_inst/edb_user_dr [59]), 
            .I1(\edb_top_inst/la0/n1814 [14]), .I2(\edb_top_inst/n1455 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3140 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3141  (.I0(\edb_top_inst/la0/n1814 [15]), 
            .I1(\edb_top_inst/la0/address_counter [15]), .I2(\edb_top_inst/n1467 ), 
            .O(\edb_top_inst/n1511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3141 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3142  (.I0(\edb_top_inst/n1511 ), .I1(\edb_top_inst/edb_user_dr [60]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3142 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3143  (.I0(\edb_top_inst/la0/n1814 [16]), 
            .I1(\edb_top_inst/la0/n1795 [1]), .I2(\edb_top_inst/n1467 ), 
            .O(\edb_top_inst/n1512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3143 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3144  (.I0(\edb_top_inst/n1512 ), .I1(\edb_top_inst/edb_user_dr [61]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3144 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3145  (.I0(\edb_top_inst/la0/n1795 [2]), .I1(\edb_top_inst/la0/n1814 [17]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3145 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3146  (.I0(\edb_top_inst/n1513 ), .I1(\edb_top_inst/edb_user_dr [62]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3146 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3147  (.I0(\edb_top_inst/la0/n1795 [3]), .I1(\edb_top_inst/la0/n1814 [18]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3147 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3148  (.I0(\edb_top_inst/n1514 ), .I1(\edb_top_inst/edb_user_dr [63]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3148 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3149  (.I0(\edb_top_inst/la0/n1795 [4]), .I1(\edb_top_inst/la0/n1814 [19]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3149 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3150  (.I0(\edb_top_inst/n1515 ), .I1(\edb_top_inst/edb_user_dr [64]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3150 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3151  (.I0(\edb_top_inst/la0/n1795 [5]), .I1(\edb_top_inst/la0/n1814 [20]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3151 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3152  (.I0(\edb_top_inst/n1516 ), .I1(\edb_top_inst/edb_user_dr [65]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3152 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3153  (.I0(\edb_top_inst/la0/n1795 [6]), .I1(\edb_top_inst/la0/n1814 [21]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3153 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3154  (.I0(\edb_top_inst/n1517 ), .I1(\edb_top_inst/edb_user_dr [66]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3154 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3155  (.I0(\edb_top_inst/la0/n1795 [7]), .I1(\edb_top_inst/la0/n1814 [22]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3155 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3156  (.I0(\edb_top_inst/n1518 ), .I1(\edb_top_inst/edb_user_dr [67]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3156 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3157  (.I0(\edb_top_inst/la0/n1795 [8]), .I1(\edb_top_inst/la0/n1814 [23]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3157 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3158  (.I0(\edb_top_inst/n1519 ), .I1(\edb_top_inst/edb_user_dr [68]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3158 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3159  (.I0(\edb_top_inst/la0/n1795 [9]), .I1(\edb_top_inst/la0/n1814 [24]), 
            .I2(\edb_top_inst/n1467 ), .O(\edb_top_inst/n1520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3159 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3160  (.I0(\edb_top_inst/n1520 ), .I1(\edb_top_inst/edb_user_dr [69]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_addr_counter [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3160 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3175  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/n1961 [1]), 
            .O(\edb_top_inst/la0/n1975 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3175 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3176  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/n1961 [2]), 
            .O(\edb_top_inst/la0/n1975 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3176 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3177  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/n1961 [3]), 
            .O(\edb_top_inst/la0/n1975 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3177 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3178  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/n1961 [4]), 
            .O(\edb_top_inst/la0/n1975 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3178 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3179  (.I0(\edb_top_inst/n1484 ), .I1(\edb_top_inst/la0/n1961 [5]), 
            .O(\edb_top_inst/la0/n1975 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3179 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3180  (.I0(\edb_top_inst/edb_user_dr [30]), 
            .I1(\edb_top_inst/la0/word_count [1]), .I2(\edb_top_inst/la0/word_count [0]), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3180 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__3181  (.I0(\edb_top_inst/la0/word_count [0]), 
            .I1(\edb_top_inst/la0/word_count [1]), .O(\edb_top_inst/n1528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3181 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3182  (.I0(\edb_top_inst/edb_user_dr [31]), 
            .I1(\edb_top_inst/la0/word_count [2]), .I2(\edb_top_inst/n1528 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3182 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3183  (.I0(\edb_top_inst/la0/word_count [2]), 
            .I1(\edb_top_inst/n1528 ), .I2(\edb_top_inst/la0/word_count [3]), 
            .O(\edb_top_inst/n1529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3183 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3184  (.I0(\edb_top_inst/n1529 ), .I1(\edb_top_inst/edb_user_dr [32]), 
            .I2(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3184 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3185  (.I0(\edb_top_inst/edb_user_dr [33]), 
            .I1(\edb_top_inst/la0/word_count [4]), .I2(\edb_top_inst/n1436 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3185 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3186  (.I0(\edb_top_inst/la0/word_count [4]), 
            .I1(\edb_top_inst/n1436 ), .O(\edb_top_inst/n1530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3186 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3187  (.I0(\edb_top_inst/edb_user_dr [34]), 
            .I1(\edb_top_inst/la0/word_count [5]), .I2(\edb_top_inst/n1530 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3187 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3188  (.I0(\edb_top_inst/la0/word_count [5]), 
            .I1(\edb_top_inst/n1530 ), .O(\edb_top_inst/n1531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3188 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3189  (.I0(\edb_top_inst/edb_user_dr [35]), 
            .I1(\edb_top_inst/la0/word_count [6]), .I2(\edb_top_inst/n1531 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3189 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3190  (.I0(\edb_top_inst/la0/word_count [6]), 
            .I1(\edb_top_inst/n1531 ), .O(\edb_top_inst/n1532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3190 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3191  (.I0(\edb_top_inst/edb_user_dr [36]), 
            .I1(\edb_top_inst/la0/word_count [7]), .I2(\edb_top_inst/n1532 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3191 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3192  (.I0(\edb_top_inst/n1435 ), .I1(\edb_top_inst/n1436 ), 
            .O(\edb_top_inst/n1533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3192 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3193  (.I0(\edb_top_inst/edb_user_dr [37]), 
            .I1(\edb_top_inst/la0/word_count [8]), .I2(\edb_top_inst/n1533 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3193 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3194  (.I0(\edb_top_inst/la0/word_count [8]), 
            .I1(\edb_top_inst/n1533 ), .O(\edb_top_inst/n1534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3194 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3195  (.I0(\edb_top_inst/edb_user_dr [38]), 
            .I1(\edb_top_inst/la0/word_count [9]), .I2(\edb_top_inst/n1534 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3195 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3196  (.I0(\edb_top_inst/la0/word_count [9]), 
            .I1(\edb_top_inst/n1534 ), .O(\edb_top_inst/n1535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3196 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3197  (.I0(\edb_top_inst/edb_user_dr [39]), 
            .I1(\edb_top_inst/la0/word_count [10]), .I2(\edb_top_inst/n1535 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3197 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3198  (.I0(\edb_top_inst/la0/word_count [10]), 
            .I1(\edb_top_inst/n1535 ), .O(\edb_top_inst/n1536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3198 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3199  (.I0(\edb_top_inst/edb_user_dr [40]), 
            .I1(\edb_top_inst/la0/word_count [11]), .I2(\edb_top_inst/n1536 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3199 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3200  (.I0(\edb_top_inst/n1434 ), .I1(\edb_top_inst/n1533 ), 
            .O(\edb_top_inst/n1537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3200 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3201  (.I0(\edb_top_inst/edb_user_dr [41]), 
            .I1(\edb_top_inst/la0/word_count [12]), .I2(\edb_top_inst/n1537 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3201 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3202  (.I0(\edb_top_inst/la0/word_count [12]), 
            .I1(\edb_top_inst/n1537 ), .O(\edb_top_inst/n1538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3202 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3203  (.I0(\edb_top_inst/edb_user_dr [42]), 
            .I1(\edb_top_inst/la0/word_count [13]), .I2(\edb_top_inst/n1538 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3203 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3204  (.I0(\edb_top_inst/la0/word_count [13]), 
            .I1(\edb_top_inst/n1538 ), .O(\edb_top_inst/n1539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3204 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3205  (.I0(\edb_top_inst/edb_user_dr [43]), 
            .I1(\edb_top_inst/la0/word_count [14]), .I2(\edb_top_inst/n1539 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3205 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3206  (.I0(\edb_top_inst/la0/word_count [14]), 
            .I1(\edb_top_inst/n1539 ), .O(\edb_top_inst/n1540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3206 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3207  (.I0(\edb_top_inst/edb_user_dr [44]), 
            .I1(\edb_top_inst/la0/word_count [15]), .I2(\edb_top_inst/n1540 ), 
            .I3(\edb_top_inst/n1455 ), .O(\edb_top_inst/la0/data_to_word_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3207 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3208  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n1541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3208 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__3209  (.I0(\edb_top_inst/n1541 ), .I1(\edb_top_inst/la0/la_trig_mask [1]), 
            .I2(\edb_top_inst/la0/internal_register_select [0]), .I3(\edb_top_inst/n1498 ), 
            .O(\edb_top_inst/n1542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3209 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3211  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3211 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3212  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [1]), 
            .I2(\edb_top_inst/n1542 ), .I3(\edb_top_inst/n1544 ), .O(\edb_top_inst/n1545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3212 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3213  (.I0(\edb_top_inst/n1545 ), .I1(\edb_top_inst/la0/data_from_biu [1]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3213 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__3214  (.I0(\edb_top_inst/n1546 ), .I1(\edb_top_inst/la0/data_out_shift_reg [2]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3214 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3215  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n1547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3215 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3216  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [2]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3216 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3217  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n1547 ), .I2(\edb_top_inst/n1498 ), .I3(\edb_top_inst/n1548 ), 
            .O(\edb_top_inst/n1549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3217 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3218  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3218 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3219  (.I0(\edb_top_inst/la0/la_trig_mask [2]), 
            .I1(\edb_top_inst/n1550 ), .O(\edb_top_inst/n1551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3219 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3220  (.I0(\edb_top_inst/n1551 ), .I1(\edb_top_inst/n1549 ), 
            .I2(\edb_top_inst/la0/data_from_biu [2]), .I3(\edb_top_inst/n1505 ), 
            .O(\edb_top_inst/n1552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3220 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__3221  (.I0(\edb_top_inst/n1552 ), .I1(\edb_top_inst/la0/data_out_shift_reg [3]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3221 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3222  (.I0(\edb_top_inst/la0/skip_count [3]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3222 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3223  (.I0(\edb_top_inst/la0/la_sample_cnt [0]), 
            .I1(\edb_top_inst/la0/la_trig_mask [3]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3223 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3224  (.I0(\edb_top_inst/n1554 ), .I1(\edb_top_inst/n1553 ), 
            .I2(\edb_top_inst/la0/data_from_biu [3]), .I3(\edb_top_inst/n1505 ), 
            .O(\edb_top_inst/n1555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3224 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__3225  (.I0(\edb_top_inst/n1555 ), .I1(\edb_top_inst/la0/data_out_shift_reg [4]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3225 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3226  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [4]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3226 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3227  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [4]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1556 ), .O(\edb_top_inst/n1557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3227 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3228  (.I0(\edb_top_inst/n1557 ), .I1(\edb_top_inst/la0/data_from_biu [4]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3228 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__3229  (.I0(\edb_top_inst/n1558 ), .I1(\edb_top_inst/la0/data_out_shift_reg [5]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3229 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3230  (.I0(\edb_top_inst/la0/skip_count [5]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3230 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3231  (.I0(\edb_top_inst/la0/la_sample_cnt [2]), 
            .I1(\edb_top_inst/la0/la_trig_mask [5]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3231 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3232  (.I0(\edb_top_inst/n1560 ), .I1(\edb_top_inst/n1559 ), 
            .I2(\edb_top_inst/la0/data_from_biu [5]), .I3(\edb_top_inst/n1505 ), 
            .O(\edb_top_inst/n1561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3232 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__3233  (.I0(\edb_top_inst/n1561 ), .I1(\edb_top_inst/la0/data_out_shift_reg [6]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3233 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3234  (.I0(\edb_top_inst/la0/la_sample_cnt [3]), 
            .I1(\edb_top_inst/la0/la_trig_mask [6]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .O(\edb_top_inst/n1562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3234 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3235  (.I0(\edb_top_inst/la0/skip_count [6]), 
            .I1(\edb_top_inst/n1501 ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3235 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__3236  (.I0(\edb_top_inst/n1563 ), .I1(\edb_top_inst/n1562 ), 
            .I2(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3236 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3237  (.I0(\edb_top_inst/n1564 ), .I1(\edb_top_inst/la0/data_from_biu [6]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3237 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3238  (.I0(\edb_top_inst/n1565 ), .I1(\edb_top_inst/la0/data_out_shift_reg [7]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3238 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3239  (.I0(\edb_top_inst/la0/skip_count [7]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3239 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3240  (.I0(\edb_top_inst/la0/la_sample_cnt [4]), 
            .I1(\edb_top_inst/la0/la_trig_mask [7]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .O(\edb_top_inst/n1567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3240 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3241  (.I0(\edb_top_inst/n1503 ), .I1(\edb_top_inst/n1566 ), 
            .I2(\edb_top_inst/n1567 ), .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3241 .LUTMASK = 16'h0fee;
    EFX_LUT4 \edb_top_inst/LUT__3242  (.I0(\edb_top_inst/n1568 ), .I1(\edb_top_inst/la0/data_from_biu [7]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3242 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3243  (.I0(\edb_top_inst/n1569 ), .I1(\edb_top_inst/la0/data_out_shift_reg [8]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3243 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3244  (.I0(\edb_top_inst/la0/la_sample_cnt [5]), 
            .I1(\edb_top_inst/la0/la_trig_mask [8]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .O(\edb_top_inst/n1570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3244 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3245  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/n1501 ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3245 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__3246  (.I0(\edb_top_inst/n1571 ), .I1(\edb_top_inst/n1570 ), 
            .I2(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3246 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3247  (.I0(\edb_top_inst/n1572 ), .I1(\edb_top_inst/la0/data_from_biu [8]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3247 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3248  (.I0(\edb_top_inst/n1573 ), .I1(\edb_top_inst/la0/data_out_shift_reg [9]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3248 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3249  (.I0(\edb_top_inst/la0/la_sample_cnt [6]), 
            .I1(\edb_top_inst/la0/la_trig_mask [9]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .O(\edb_top_inst/n1574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3249 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3250  (.I0(\edb_top_inst/la0/skip_count [9]), 
            .I1(\edb_top_inst/n1501 ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3250 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__3251  (.I0(\edb_top_inst/n1575 ), .I1(\edb_top_inst/n1574 ), 
            .I2(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3251 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3252  (.I0(\edb_top_inst/n1576 ), .I1(\edb_top_inst/la0/data_from_biu [9]), 
            .I2(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3252 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__3253  (.I0(\edb_top_inst/n1577 ), .I1(\edb_top_inst/la0/data_out_shift_reg [10]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3253 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3254  (.I0(\edb_top_inst/la0/la_sample_cnt [7]), 
            .I1(\edb_top_inst/la0/la_trig_mask [10]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3254 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3255  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [10]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1578 ), .O(\edb_top_inst/n1579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3255 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3256  (.I0(\edb_top_inst/n1579 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [11]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3256 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3257  (.I0(\edb_top_inst/la0/la_sample_cnt [8]), 
            .I1(\edb_top_inst/la0/la_trig_mask [11]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3257 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3258  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [11]), 
            .I2(\edb_top_inst/n1580 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3258 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3259  (.I0(\edb_top_inst/n1581 ), .I1(\edb_top_inst/la0/data_out_shift_reg [12]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3259 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3260  (.I0(\edb_top_inst/la0/la_sample_cnt [9]), 
            .I1(\edb_top_inst/la0/la_trig_mask [12]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3260 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3261  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [12]), 
            .I2(\edb_top_inst/n1582 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3261 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3262  (.I0(\edb_top_inst/n1583 ), .I1(\edb_top_inst/la0/data_out_shift_reg [13]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3262 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3263  (.I0(\edb_top_inst/la0/la_sample_cnt [10]), 
            .I1(\edb_top_inst/la0/la_trig_mask [13]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3263 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3264  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [13]), 
            .I2(\edb_top_inst/n1584 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3264 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3265  (.I0(\edb_top_inst/n1585 ), .I1(\edb_top_inst/la0/data_out_shift_reg [14]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3265 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3266  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [14]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3266 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3267  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [14]), 
            .I2(\edb_top_inst/n1586 ), .O(\edb_top_inst/n1587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3267 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3268  (.I0(\edb_top_inst/n1587 ), .I1(\edb_top_inst/la0/data_out_shift_reg [15]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3268 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3269  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [15]), 
            .I2(\edb_top_inst/la0/la_trig_mask [15]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3269 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3270  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [16]), 
            .I2(\edb_top_inst/n1588 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3270 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3271  (.I0(\edb_top_inst/la0/skip_count [16]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3271 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3272  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [16]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1589 ), .O(\edb_top_inst/n1590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3272 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3273  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [17]), 
            .I2(\edb_top_inst/n1590 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3273 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3274  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [17]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3274 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3275  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [17]), 
            .I2(\edb_top_inst/n1591 ), .O(\edb_top_inst/n1592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3275 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3276  (.I0(\edb_top_inst/n1592 ), .I1(\edb_top_inst/la0/data_out_shift_reg [18]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3276 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3277  (.I0(\edb_top_inst/la0/skip_count [18]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3277 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3278  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [18]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1593 ), .O(\edb_top_inst/n1594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3278 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3279  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [19]), 
            .I2(\edb_top_inst/n1594 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3279 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3280  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [19]), 
            .I2(\edb_top_inst/la0/la_trig_mask [19]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3280 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3281  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [20]), 
            .I2(\edb_top_inst/n1595 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3281 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3282  (.I0(\edb_top_inst/la0/la_trig_mask [20]), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3282 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__3283  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [20]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1596 ), .O(\edb_top_inst/n1597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3283 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3284  (.I0(\edb_top_inst/n1597 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [21]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3284 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3285  (.I0(\edb_top_inst/la0/la_trig_mask [21]), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3285 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__3286  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [21]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1598 ), .O(\edb_top_inst/n1599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3286 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3287  (.I0(\edb_top_inst/n1599 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [22]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3287 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3288  (.I0(\edb_top_inst/la0/la_trig_mask [22]), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3288 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__3289  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [22]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1600 ), .O(\edb_top_inst/n1601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3289 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3290  (.I0(\edb_top_inst/n1601 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [23]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3290 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3291  (.I0(\edb_top_inst/la0/internal_register_select [0]), 
            .I1(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3291 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3293  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [23]), 
            .I2(\edb_top_inst/la0/la_trig_mask [23]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3293 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3294  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_trig_pos [0]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1604 ), .O(\edb_top_inst/n1605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3294 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3295  (.I0(\edb_top_inst/n1605 ), .I1(\edb_top_inst/la0/data_out_shift_reg [24]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3295 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3296  (.I0(\edb_top_inst/la0/la_trig_pos [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [24]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3296 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3297  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [24]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1606 ), .O(\edb_top_inst/n1607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3297 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3298  (.I0(\edb_top_inst/n1607 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [25]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3298 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3299  (.I0(\edb_top_inst/la0/la_trig_pos [2]), 
            .I1(\edb_top_inst/la0/la_trig_mask [25]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3299 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3300  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [25]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1608 ), .O(\edb_top_inst/n1609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3300 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3301  (.I0(\edb_top_inst/n1609 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [26]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3301 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3302  (.I0(\edb_top_inst/la0/la_trig_pos [3]), 
            .I1(\edb_top_inst/la0/la_trig_mask [26]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3302 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3303  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [26]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1610 ), .O(\edb_top_inst/n1611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3303 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3304  (.I0(\edb_top_inst/n1611 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [27]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3304 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3305  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [27]), 
            .I2(\edb_top_inst/la0/la_trig_mask [27]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3305 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3306  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_trig_pos [4]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1612 ), .O(\edb_top_inst/n1613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3306 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3307  (.I0(\edb_top_inst/n1613 ), .I1(\edb_top_inst/la0/data_out_shift_reg [28]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3307 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3308  (.I0(\edb_top_inst/la0/la_trig_pos [5]), 
            .I1(\edb_top_inst/la0/la_trig_mask [28]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3308 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3309  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [28]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1614 ), .O(\edb_top_inst/n1615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3309 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3310  (.I0(\edb_top_inst/n1615 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [29]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3310 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3311  (.I0(\edb_top_inst/la0/la_trig_pos [6]), 
            .I1(\edb_top_inst/la0/la_trig_mask [29]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3311 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3312  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [29]), 
            .I2(\edb_top_inst/n1616 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3312 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3313  (.I0(\edb_top_inst/n1617 ), .I1(\edb_top_inst/la0/data_out_shift_reg [30]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3313 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3314  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [30]), 
            .I2(\edb_top_inst/la0/la_trig_mask [30]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3314 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3315  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_trig_pos [7]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1618 ), .O(\edb_top_inst/n1619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3315 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3316  (.I0(\edb_top_inst/n1619 ), .I1(\edb_top_inst/la0/data_out_shift_reg [31]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3316 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3317  (.I0(\edb_top_inst/la0/la_trig_pos [8]), 
            .I1(\edb_top_inst/la0/la_trig_mask [31]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3317 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3318  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [31]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1620 ), .O(\edb_top_inst/n1621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3318 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3319  (.I0(\edb_top_inst/n1621 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [32]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3319 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3320  (.I0(\edb_top_inst/la0/la_trig_pos [9]), 
            .I1(\edb_top_inst/la0/la_trig_mask [32]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3320 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3321  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [32]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1622 ), .O(\edb_top_inst/n1623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3321 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3322  (.I0(\edb_top_inst/n1623 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [33]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3322 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3323  (.I0(\edb_top_inst/la0/la_trig_pos [10]), 
            .I1(\edb_top_inst/la0/la_trig_mask [33]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3323 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3324  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [33]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1624 ), .O(\edb_top_inst/n1625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3324 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3325  (.I0(\edb_top_inst/n1625 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [34]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3325 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3326  (.I0(\edb_top_inst/la0/la_trig_pos [11]), 
            .I1(\edb_top_inst/la0/la_trig_mask [34]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3326 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3327  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [34]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1626 ), .O(\edb_top_inst/n1627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3327 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3328  (.I0(\edb_top_inst/n1627 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [35]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3328 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3329  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [35]), 
            .I2(\edb_top_inst/la0/la_trig_mask [35]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3329 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3330  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_trig_pos [12]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1628 ), .O(\edb_top_inst/n1629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3330 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3331  (.I0(\edb_top_inst/n1629 ), .I1(\edb_top_inst/la0/data_out_shift_reg [36]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3331 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3332  (.I0(\edb_top_inst/la0/la_trig_pos [13]), 
            .I1(\edb_top_inst/la0/la_trig_mask [36]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3332 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3333  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [36]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1630 ), .O(\edb_top_inst/n1631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3333 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3334  (.I0(\edb_top_inst/n1631 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [37]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3334 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3335  (.I0(\edb_top_inst/la0/la_trig_pos [14]), 
            .I1(\edb_top_inst/la0/la_trig_mask [37]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3335 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3336  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [37]), 
            .I2(\edb_top_inst/n1502 ), .I3(\edb_top_inst/n1632 ), .O(\edb_top_inst/n1633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3336 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3337  (.I0(\edb_top_inst/n1633 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [38]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3337 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3338  (.I0(\edb_top_inst/la0/la_trig_pos [15]), 
            .I1(\edb_top_inst/la0/la_trig_mask [38]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3338 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3339  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [38]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1634 ), .O(\edb_top_inst/n1635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3339 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3340  (.I0(\edb_top_inst/n1635 ), .I1(\edb_top_inst/n1505 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg [39]), .I3(\edb_top_inst/n1508 ), 
            .O(\edb_top_inst/la0/n2194 [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3340 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3341  (.I0(\edb_top_inst/la0/la_trig_pos [16]), 
            .I1(\edb_top_inst/la0/la_trig_mask [39]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3341 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3342  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [39]), 
            .I2(\edb_top_inst/n1636 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3342 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3343  (.I0(\edb_top_inst/n1637 ), .I1(\edb_top_inst/la0/data_out_shift_reg [40]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3343 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3344  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [40]), 
            .I2(\edb_top_inst/la0/la_trig_mask [40]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3344 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3345  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_trig_pattern [0]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1638 ), .O(\edb_top_inst/n1639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3345 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3346  (.I0(\edb_top_inst/n1639 ), .I1(\edb_top_inst/la0/data_out_shift_reg [41]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3346 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3347  (.I0(\edb_top_inst/la0/la_trig_mask [41]), 
            .I1(\edb_top_inst/la0/la_trig_pattern [1]), .I2(\edb_top_inst/la0/internal_register_select [0]), 
            .I3(\edb_top_inst/n1498 ), .O(\edb_top_inst/n1640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3347 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__3348  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [41]), 
            .I2(\edb_top_inst/n1640 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/n1641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3348 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3349  (.I0(\edb_top_inst/n1641 ), .I1(\edb_top_inst/la0/data_out_shift_reg [42]), 
            .I2(\edb_top_inst/n1508 ), .O(\edb_top_inst/la0/n2194 [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3349 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3350  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [42]), 
            .I2(\edb_top_inst/la0/la_trig_mask [42]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3350 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3351  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_capture_pattern [0]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1642 ), .O(\edb_top_inst/n1643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3351 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3352  (.I0(\edb_top_inst/n1643 ), .I1(\edb_top_inst/la0/data_out_shift_reg [43]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3352 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3353  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [43]), 
            .I2(\edb_top_inst/la0/la_trig_mask [43]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3353 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3354  (.I0(\edb_top_inst/n1602 ), .I1(\edb_top_inst/la0/la_capture_pattern [1]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1644 ), .O(\edb_top_inst/n1645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3354 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3355  (.I0(\edb_top_inst/n1645 ), .I1(\edb_top_inst/la0/data_out_shift_reg [44]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3355 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3356  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3356 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3357  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [44]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1646 ), .O(\edb_top_inst/n1647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3357 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3358  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [45]), 
            .I2(\edb_top_inst/n1647 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3358 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3359  (.I0(\edb_top_inst/la0/skip_count [45]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3359 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3360  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [45]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1648 ), .O(\edb_top_inst/n1649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3360 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3361  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [46]), 
            .I2(\edb_top_inst/n1649 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3361 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3363  (.I0(\edb_top_inst/la0/skip_count [46]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3363 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3364  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [46]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1651 ), .O(\edb_top_inst/n1652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3364 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3365  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [47]), 
            .I2(\edb_top_inst/n1652 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3365 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3366  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [47]), 
            .I2(\edb_top_inst/la0/la_trig_mask [47]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3366 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3367  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [48]), 
            .I2(\edb_top_inst/n1653 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3367 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3368  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [48]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3368 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3369  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [48]), 
            .I2(\edb_top_inst/n1654 ), .O(\edb_top_inst/n1655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3369 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3370  (.I0(\edb_top_inst/n1655 ), .I1(\edb_top_inst/la0/data_out_shift_reg [49]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3370 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3371  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [49]), 
            .I2(\edb_top_inst/la0/la_trig_mask [49]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3371 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3372  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [50]), 
            .I2(\edb_top_inst/n1656 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3372 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3373  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [50]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3373 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3374  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [50]), 
            .I2(\edb_top_inst/n1657 ), .O(\edb_top_inst/n1658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3374 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3375  (.I0(\edb_top_inst/n1658 ), .I1(\edb_top_inst/la0/data_out_shift_reg [51]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3375 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3376  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [51]), 
            .I2(\edb_top_inst/la0/la_trig_mask [51]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3376 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3377  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [52]), 
            .I2(\edb_top_inst/n1659 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3377 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3378  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3378 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3379  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [52]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1660 ), .O(\edb_top_inst/n1661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3379 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3380  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [53]), 
            .I2(\edb_top_inst/n1661 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3380 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3381  (.I0(\edb_top_inst/la0/skip_count [53]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3381 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3382  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [53]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1662 ), .O(\edb_top_inst/n1663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3382 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3383  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [54]), 
            .I2(\edb_top_inst/n1663 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3383 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3384  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [54]), 
            .I2(\edb_top_inst/la0/la_trig_mask [54]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3384 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3385  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [55]), 
            .I2(\edb_top_inst/n1664 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3385 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3386  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3386 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3387  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [55]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1665 ), .O(\edb_top_inst/n1666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3387 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3388  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [56]), 
            .I2(\edb_top_inst/n1666 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3388 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3389  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [56]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3389 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3390  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [56]), 
            .I2(\edb_top_inst/n1667 ), .O(\edb_top_inst/n1668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3390 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3391  (.I0(\edb_top_inst/n1668 ), .I1(\edb_top_inst/la0/data_out_shift_reg [57]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3391 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3392  (.I0(\edb_top_inst/la0/skip_count [57]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3392 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3393  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [57]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1669 ), .O(\edb_top_inst/n1670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3393 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3394  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [58]), 
            .I2(\edb_top_inst/n1670 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3394 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3395  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3395 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3396  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [58]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1671 ), .O(\edb_top_inst/n1672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3396 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3397  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [59]), 
            .I2(\edb_top_inst/n1672 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3397 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3398  (.I0(\edb_top_inst/la0/skip_count [59]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3398 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3399  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [59]), 
            .I2(\edb_top_inst/n1544 ), .I3(\edb_top_inst/n1673 ), .O(\edb_top_inst/n1674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3399 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3400  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [60]), 
            .I2(\edb_top_inst/n1674 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3400 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3401  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [60]), 
            .I2(\edb_top_inst/n1502 ), .O(\edb_top_inst/n1675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3401 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3402  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [60]), 
            .I2(\edb_top_inst/n1675 ), .O(\edb_top_inst/n1676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3402 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3403  (.I0(\edb_top_inst/n1676 ), .I1(\edb_top_inst/la0/data_out_shift_reg [61]), 
            .I2(\edb_top_inst/n1507 ), .I3(\edb_top_inst/n1505 ), .O(\edb_top_inst/la0/n2194 [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3403 .LUTMASK = 16'h5c00;
    EFX_LUT4 \edb_top_inst/LUT__3404  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [61]), 
            .I2(\edb_top_inst/la0/la_trig_mask [61]), .I3(\edb_top_inst/n1550 ), 
            .O(\edb_top_inst/n1677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3404 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3405  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [62]), 
            .I2(\edb_top_inst/n1677 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3405 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3406  (.I0(\edb_top_inst/la0/skip_count [62]), 
            .I1(\edb_top_inst/n1501 ), .O(\edb_top_inst/n1678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3406 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3407  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [62]), 
            .I2(\edb_top_inst/n1503 ), .I3(\edb_top_inst/n1678 ), .O(\edb_top_inst/n1679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3407 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3408  (.I0(\edb_top_inst/n1505 ), .I1(\edb_top_inst/la0/data_out_shift_reg [63]), 
            .I2(\edb_top_inst/n1679 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3408 .LUTMASK = 16'h0f88;
    EFX_LUT4 \edb_top_inst/LUT__3409  (.I0(\edb_top_inst/n1501 ), .I1(\edb_top_inst/la0/skip_count [63]), 
            .I2(\edb_top_inst/n1544 ), .O(\edb_top_inst/n1680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3409 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3410  (.I0(\edb_top_inst/n1550 ), .I1(\edb_top_inst/la0/la_trig_mask [63]), 
            .I2(\edb_top_inst/n1680 ), .I3(\edb_top_inst/n1507 ), .O(\edb_top_inst/la0/n2194 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3410 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3411  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n1441 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/la0/module_state [1]), 
            .O(\edb_top_inst/n1681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3411 .LUTMASK = 16'hf077;
    EFX_LUT4 \edb_top_inst/LUT__3412  (.I0(\edb_top_inst/n1442 ), .I1(\edb_top_inst/n1429 ), 
            .O(\edb_top_inst/n1682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3412 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3413  (.I0(\edb_top_inst/n1682 ), .I1(\edb_top_inst/n1681 ), 
            .I2(\edb_top_inst/la0/module_state [3]), .I3(\edb_top_inst/la0/module_state [2]), 
            .O(\edb_top_inst/n1683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3413 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3414  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n1450 ), 
            .O(\edb_top_inst/n1684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3414 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3415  (.I0(\edb_top_inst/n1438 ), .I1(\edb_top_inst/n1683 ), 
            .I2(\edb_top_inst/n1684 ), .I3(\edb_top_inst/la0/module_state [0]), 
            .O(\edb_top_inst/n1685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3415 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__3416  (.I0(\edb_top_inst/n1684 ), .I1(\edb_top_inst/n1683 ), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/n1685 ), 
            .O(\edb_top_inst/la0/module_next_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3416 .LUTMASK = 16'he0ff;
    EFX_LUT4 \edb_top_inst/LUT__3417  (.I0(\edb_top_inst/la0/module_state [0]), 
            .I1(\edb_top_inst/n1485 ), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(jtag_inst1_UPDATE), .O(\edb_top_inst/n1686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3417 .LUTMASK = 16'h0071;
    EFX_LUT4 \edb_top_inst/LUT__3418  (.I0(\edb_top_inst/n1438 ), .I1(\edb_top_inst/n1445 ), 
            .I2(\edb_top_inst/n1684 ), .I3(\edb_top_inst/n1479 ), .O(\edb_top_inst/n1687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3418 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__3419  (.I0(\edb_top_inst/n1478 ), .I1(\edb_top_inst/n1686 ), 
            .I2(\edb_top_inst/n1687 ), .I3(\edb_top_inst/n1489 ), .O(\edb_top_inst/la0/module_next_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3419 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__3420  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n1438 ), 
            .I2(\edb_top_inst/n1476 ), .I3(\edb_top_inst/n1489 ), .O(\edb_top_inst/n1688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3420 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3421  (.I0(\edb_top_inst/n1438 ), .I1(\edb_top_inst/n1445 ), 
            .I2(\edb_top_inst/n1684 ), .I3(\edb_top_inst/n1688 ), .O(\edb_top_inst/la0/module_next_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3421 .LUTMASK = 16'hffb0;
    EFX_LUT4 \edb_top_inst/LUT__3422  (.I0(\edb_top_inst/la0/crc_data_out [1]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3422 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3423  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/n1450 ), 
            .O(\edb_top_inst/n1689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3423 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3424  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n1490 ), .I2(\edb_top_inst/n1689 ), .O(\edb_top_inst/ceg_net11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3424 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3425  (.I0(\edb_top_inst/la0/crc_data_out [2]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3425 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3426  (.I0(\edb_top_inst/la0/crc_data_out [3]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3426 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3427  (.I0(\edb_top_inst/la0/crc_data_out [4]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3427 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3428  (.I0(\edb_top_inst/la0/crc_data_out [5]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3428 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3429  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg [0]), 
            .I2(\edb_top_inst/la0/module_state [1]), .I3(\edb_top_inst/la0/crc_data_out [0]), 
            .O(\edb_top_inst/n1690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3429 .LUTMASK = 16'hac53;
    EFX_LUT4 \edb_top_inst/LUT__3430  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/n1690 ), 
            .I3(\edb_top_inst/n1489 ), .O(\edb_top_inst/n1691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3430 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__3431  (.I0(\edb_top_inst/la0/module_next_state [0]), 
            .I1(\edb_top_inst/la0/module_state [0]), .I2(\edb_top_inst/la0/module_state [1]), 
            .I3(\edb_top_inst/n1691 ), .O(\edb_top_inst/n1692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3431 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__3432  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [6]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3432 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3433  (.I0(\edb_top_inst/la0/crc_data_out [7]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3433 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3434  (.I0(\edb_top_inst/la0/crc_data_out [8]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3434 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3435  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [9]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3435 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3436  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [10]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3436 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3437  (.I0(\edb_top_inst/la0/crc_data_out [11]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3437 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3438  (.I0(\edb_top_inst/la0/crc_data_out [12]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3438 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3439  (.I0(\edb_top_inst/la0/crc_data_out [13]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3439 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3440  (.I0(\edb_top_inst/la0/crc_data_out [14]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3440 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3441  (.I0(\edb_top_inst/la0/crc_data_out [15]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3441 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3442  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [16]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3442 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3443  (.I0(\edb_top_inst/la0/crc_data_out [17]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3443 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3444  (.I0(\edb_top_inst/la0/crc_data_out [18]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3444 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3445  (.I0(\edb_top_inst/la0/crc_data_out [19]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3445 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3446  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [20]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3446 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3447  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [21]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3447 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3448  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [22]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3448 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3449  (.I0(\edb_top_inst/la0/crc_data_out [23]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3449 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3450  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [24]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3450 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3451  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [25]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3451 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3452  (.I0(\edb_top_inst/la0/crc_data_out [26]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3452 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3453  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [27]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3453 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3454  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [28]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3454 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3455  (.I0(\edb_top_inst/la0/crc_data_out [29]), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n118 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3455 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3456  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [30]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3456 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3457  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out [31]), .I2(\edb_top_inst/n1692 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n118 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3457 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3458  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n1692 ), .O(\edb_top_inst/la0/axi_crc_i/n118 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3458 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3459  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3459 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3460  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3460 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3461  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3461 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__3462  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3462 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3463  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n1693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3463 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__3464  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/n1693 ), .O(\edb_top_inst/n1694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3464 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__3465  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/n1695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3465 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__3466  (.I0(\edb_top_inst/n1695 ), .I1(\edb_top_inst/n1694 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3466 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3467  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3467 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3468  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [0]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3468 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3469  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), .O(\edb_top_inst/n1696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3469 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__3470  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/n1696 ), .O(\edb_top_inst/n1697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3470 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__3471  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I2(\edb_top_inst/n1697 ), .O(\edb_top_inst/n1698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3471 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__3472  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I2(\edb_top_inst/n1698 ), .O(\edb_top_inst/n1699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3472 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__3473  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/n1699 ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/n1700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3473 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__3474  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I2(\edb_top_inst/n1700 ), .O(\edb_top_inst/n1701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3474 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__3475  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I2(\edb_top_inst/n1701 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3475 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__3476  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/n1702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3476 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3477  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/n1703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3477 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3478  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/n1704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3478 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3479  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/n1705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3479 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3480  (.I0(\edb_top_inst/n1702 ), .I1(\edb_top_inst/n1703 ), 
            .I2(\edb_top_inst/n1704 ), .I3(\edb_top_inst/n1705 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3480 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__3481  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n1706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3481 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__3482  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n1707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3482 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3483  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [0]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [0]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [1]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [1]), 
            .O(\edb_top_inst/n1708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3483 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3484  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [4]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [5]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [5]), 
            .O(\edb_top_inst/n1709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3484 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3485  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [6]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [7]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [7]), 
            .O(\edb_top_inst/n1710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3485 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3486  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [2]), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2 [3]), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 [3]), 
            .O(\edb_top_inst/n1711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3486 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3487  (.I0(\edb_top_inst/n1708 ), .I1(\edb_top_inst/n1709 ), 
            .I2(\edb_top_inst/n1710 ), .I3(\edb_top_inst/n1711 ), .O(\edb_top_inst/n1712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3487 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3488  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/n1707 ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [0]), 
            .I3(\edb_top_inst/n1712 ), .O(\edb_top_inst/n1713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2f75, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3488 .LUTMASK = 16'h2f75;
    EFX_LUT4 \edb_top_inst/LUT__3489  (.I0(\edb_top_inst/n1713 ), .I1(\edb_top_inst/n1706 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3489 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3490  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3490 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3491  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3491 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3492  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3492 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3493  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3493 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3494  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3494 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3495  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3495 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3496  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n32 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3496 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3497  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [1]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3497 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3498  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [2]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [2]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3498 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3499  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [3]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [3]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3499 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3500  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [4]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [4]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3500 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3501  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [5]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [5]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3501 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3502  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [6]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [6]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3502 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3503  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1 [7]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr [7]), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n14 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3503 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3504  (.I0(\edb_top_inst/la0/la_trig_mask [1]), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask [0]), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n1714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3504 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3505  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask [1]), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask [0]), .O(\edb_top_inst/n1715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3505 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__3506  (.I0(\edb_top_inst/n1714 ), .I1(\edb_top_inst/n1715 ), 
            .I2(\edb_top_inst/la0/la_trig_pattern [0]), .I3(\edb_top_inst/la0/la_trig_pattern [1]), 
            .O(\edb_top_inst/n1716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ca3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3506 .LUTMASK = 16'h5ca3;
    EFX_LUT4 \edb_top_inst/LUT__3507  (.I0(\edb_top_inst/la0/la_trig_mask [1]), 
            .I1(\edb_top_inst/la0/la_trig_mask [0]), .I2(\edb_top_inst/n1716 ), 
            .O(\edb_top_inst/la0/trigger_tu/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3507 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__3508  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .I2(\edb_top_inst/la0/skip_count [2]), 
            .I3(\edb_top_inst/la0/skip_count [3]), .O(\edb_top_inst/n1717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3508 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3509  (.I0(\edb_top_inst/la0/skip_count [4]), 
            .I1(\edb_top_inst/la0/skip_count [5]), .I2(\edb_top_inst/la0/skip_count [6]), 
            .I3(\edb_top_inst/la0/skip_count [7]), .O(\edb_top_inst/n1718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3509 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3510  (.I0(\edb_top_inst/la0/skip_count [9]), 
            .I1(\edb_top_inst/la0/skip_count [10]), .I2(\edb_top_inst/la0/skip_count [11]), 
            .I3(\edb_top_inst/la0/skip_count [12]), .O(\edb_top_inst/n1719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3510 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3511  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/n1717 ), .I2(\edb_top_inst/n1718 ), .I3(\edb_top_inst/n1719 ), 
            .O(\edb_top_inst/n1720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3511 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3512  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/la0/skip_count [14]), .I2(\edb_top_inst/la0/skip_count [15]), 
            .I3(\edb_top_inst/la0/skip_count [16]), .O(\edb_top_inst/n1721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3512 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3513  (.I0(\edb_top_inst/la0/skip_count [18]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18]), 
            .O(\edb_top_inst/n1722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3513 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3514  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/n1720 ), .I2(\edb_top_inst/n1721 ), .I3(\edb_top_inst/n1722 ), 
            .O(\edb_top_inst/n1723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3514 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3515  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/la0/skip_count [18]), .I2(\edb_top_inst/la0/skip_count [19]), 
            .I3(\edb_top_inst/la0/skip_count [20]), .O(\edb_top_inst/n1724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3515 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3516  (.I0(\edb_top_inst/la0/skip_count [21]), 
            .I1(\edb_top_inst/n1721 ), .I2(\edb_top_inst/n1724 ), .O(\edb_top_inst/n1725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3516 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3517  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/skip_count [27]), .I2(\edb_top_inst/la0/skip_count [28]), 
            .I3(\edb_top_inst/la0/skip_count [29]), .O(\edb_top_inst/n1726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3517 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3518  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/skip_count [23]), .I2(\edb_top_inst/la0/skip_count [24]), 
            .I3(\edb_top_inst/la0/skip_count [25]), .O(\edb_top_inst/n1727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3518 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3519  (.I0(\edb_top_inst/la0/skip_count [30]), 
            .I1(\edb_top_inst/la0/skip_count [31]), .I2(\edb_top_inst/n1726 ), 
            .I3(\edb_top_inst/n1727 ), .O(\edb_top_inst/n1728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3519 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3520  (.I0(\edb_top_inst/la0/skip_count [38]), 
            .I1(\edb_top_inst/la0/skip_count [39]), .O(\edb_top_inst/n1729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3520 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3521  (.I0(\edb_top_inst/la0/skip_count [34]), 
            .I1(\edb_top_inst/la0/skip_count [35]), .I2(\edb_top_inst/la0/skip_count [36]), 
            .I3(\edb_top_inst/la0/skip_count [37]), .O(\edb_top_inst/n1730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3521 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3522  (.I0(\edb_top_inst/la0/skip_count [32]), 
            .I1(\edb_top_inst/la0/skip_count [33]), .I2(\edb_top_inst/n1729 ), 
            .I3(\edb_top_inst/n1730 ), .O(\edb_top_inst/n1731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3522 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3523  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1728 ), .I3(\edb_top_inst/n1731 ), .O(\edb_top_inst/n1732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3523 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3524  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/skip_count [41]), .I2(\edb_top_inst/la0/skip_count [42]), 
            .I3(\edb_top_inst/la0/skip_count [43]), .O(\edb_top_inst/n1733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3524 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3525  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1733 ), 
            .I2(\edb_top_inst/la0/skip_count [44]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .O(\edb_top_inst/n1734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3525 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3526  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/skip_count [41]), .O(\edb_top_inst/n1735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3526 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3527  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1735 ), 
            .I2(\edb_top_inst/la0/skip_count [42]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42]), 
            .O(\edb_top_inst/n1736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3527 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3528  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/la0/skip_count [45]), .I2(\edb_top_inst/la0/skip_count [46]), 
            .O(\edb_top_inst/n1737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3528 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3529  (.I0(\edb_top_inst/la0/skip_count [47]), 
            .I1(\edb_top_inst/la0/skip_count [48]), .I2(\edb_top_inst/n1733 ), 
            .I3(\edb_top_inst/n1737 ), .O(\edb_top_inst/n1738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3529 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3530  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1738 ), 
            .O(\edb_top_inst/n1739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3530 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3531  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49]), 
            .O(\edb_top_inst/n1740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3531 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3532  (.I0(\edb_top_inst/n1739 ), .I1(\edb_top_inst/n1740 ), 
            .I2(\edb_top_inst/n1734 ), .I3(\edb_top_inst/n1736 ), .O(\edb_top_inst/n1741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3532 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__3533  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/n1732 ), .I2(\edb_top_inst/la0/skip_count [41]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41]), 
            .O(\edb_top_inst/n1742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb44b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3533 .LUTMASK = 16'hb44b;
    EFX_LUT4 \edb_top_inst/LUT__3534  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/skip_count [50]), .I2(\edb_top_inst/la0/skip_count [51]), 
            .I3(\edb_top_inst/la0/skip_count [52]), .O(\edb_top_inst/n1743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3534 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3535  (.I0(\edb_top_inst/la0/skip_count [53]), 
            .I1(\edb_top_inst/n1738 ), .I2(\edb_top_inst/n1743 ), .O(\edb_top_inst/n1744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3535 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3536  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1744 ), 
            .I2(\edb_top_inst/la0/skip_count [54]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54]), 
            .O(\edb_top_inst/n1745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3536 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3537  (.I0(\edb_top_inst/n1726 ), .I1(\edb_top_inst/n1727 ), 
            .O(\edb_top_inst/n1746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3537 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3538  (.I0(\edb_top_inst/la0/skip_count [30]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30]), 
            .O(\edb_top_inst/n1747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3538 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3539  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1746 ), .I3(\edb_top_inst/n1747 ), .O(\edb_top_inst/n1748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3539 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__3540  (.I0(\edb_top_inst/la0/skip_count [32]), 
            .I1(\edb_top_inst/n1720 ), .I2(\edb_top_inst/n1725 ), .I3(\edb_top_inst/n1728 ), 
            .O(\edb_top_inst/n1749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3540 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3541  (.I0(\edb_top_inst/la0/skip_count [33]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33]), 
            .I2(\edb_top_inst/n1749 ), .I3(\edb_top_inst/n1748 ), .O(\edb_top_inst/n1750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3541 .LUTMASK = 16'h6900;
    EFX_LUT4 \edb_top_inst/LUT__3542  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .O(\edb_top_inst/n1751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3542 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3543  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/skip_count [27]), .I2(\edb_top_inst/la0/skip_count [28]), 
            .I3(\edb_top_inst/n1727 ), .O(\edb_top_inst/n1752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3543 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3544  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/n1727 ), .O(\edb_top_inst/n1753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3544 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3545  (.I0(\edb_top_inst/la0/skip_count [27]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27]), 
            .O(\edb_top_inst/n1754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3545 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3546  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1753 ), .I3(\edb_top_inst/n1754 ), .O(\edb_top_inst/n1755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3546 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__3547  (.I0(\edb_top_inst/la0/skip_count [29]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29]), 
            .O(\edb_top_inst/n1756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3547 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3548  (.I0(\edb_top_inst/n1751 ), .I1(\edb_top_inst/n1752 ), 
            .I2(\edb_top_inst/n1756 ), .I3(\edb_top_inst/n1755 ), .O(\edb_top_inst/n1757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3548 .LUTMASK = 16'h7800;
    EFX_LUT4 \edb_top_inst/LUT__3549  (.I0(\edb_top_inst/n1742 ), .I1(\edb_top_inst/n1745 ), 
            .I2(\edb_top_inst/n1750 ), .I3(\edb_top_inst/n1757 ), .O(\edb_top_inst/n1758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3549 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3550  (.I0(\edb_top_inst/la0/skip_count [10]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10]), 
            .O(\edb_top_inst/n1759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3550 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3551  (.I0(\edb_top_inst/n1717 ), .I1(\edb_top_inst/n1718 ), 
            .O(\edb_top_inst/n1760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3551 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3552  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/n1760 ), .O(\edb_top_inst/n1761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3552 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3553  (.I0(\edb_top_inst/la0/skip_count [9]), 
            .I1(\edb_top_inst/n1759 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9]), 
            .I3(\edb_top_inst/n1761 ), .O(\edb_top_inst/n1762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3553 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3554  (.I0(\edb_top_inst/la0/skip_count [34]), 
            .I1(\edb_top_inst/la0/skip_count [35]), .O(\edb_top_inst/n1763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3554 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3555  (.I0(\edb_top_inst/la0/skip_count [30]), 
            .I1(\edb_top_inst/la0/skip_count [31]), .O(\edb_top_inst/n1764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3555 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3556  (.I0(\edb_top_inst/la0/skip_count [32]), 
            .I1(\edb_top_inst/la0/skip_count [33]), .O(\edb_top_inst/n1765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3556 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3557  (.I0(\edb_top_inst/n1726 ), .I1(\edb_top_inst/n1727 ), 
            .I2(\edb_top_inst/n1764 ), .I3(\edb_top_inst/n1765 ), .O(\edb_top_inst/n1766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3557 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3558  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1766 ), .O(\edb_top_inst/n1767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3558 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3559  (.I0(\edb_top_inst/n1763 ), .I1(\edb_top_inst/n1767 ), 
            .I2(\edb_top_inst/la0/skip_count [36]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36]), 
            .O(\edb_top_inst/n1768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3559 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3560  (.I0(\edb_top_inst/la0/skip_count [40]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40]), 
            .O(\edb_top_inst/n1769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3560 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3561  (.I0(\edb_top_inst/la0/skip_count [34]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34]), 
            .O(\edb_top_inst/n1770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3561 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3562  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1770 ), 
            .I2(\edb_top_inst/n1767 ), .I3(\edb_top_inst/n1769 ), .O(\edb_top_inst/n1771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3562 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__3563  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26]), 
            .O(\edb_top_inst/n1772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3563 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3564  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1727 ), .I3(\edb_top_inst/n1772 ), .O(\edb_top_inst/n1773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3564 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__3565  (.I0(\edb_top_inst/la0/skip_count [26]), 
            .I1(\edb_top_inst/la0/skip_count [27]), .I2(\edb_top_inst/n1727 ), 
            .O(\edb_top_inst/n1774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3565 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3566  (.I0(\edb_top_inst/la0/skip_count [28]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28]), 
            .O(\edb_top_inst/n1775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3566 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3567  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1774 ), .I3(\edb_top_inst/n1775 ), .O(\edb_top_inst/n1776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3567 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__3568  (.I0(\edb_top_inst/la0/skip_count [37]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37]), 
            .O(\edb_top_inst/n1777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3568 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3569  (.I0(\edb_top_inst/la0/skip_count [36]), 
            .I1(\edb_top_inst/n1763 ), .O(\edb_top_inst/n1778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3569 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3570  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1778 ), .I3(\edb_top_inst/n1766 ), .O(\edb_top_inst/n1779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3570 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3571  (.I0(\edb_top_inst/n1777 ), .I1(\edb_top_inst/n1779 ), 
            .I2(\edb_top_inst/n1773 ), .I3(\edb_top_inst/n1776 ), .O(\edb_top_inst/n1780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3571 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__3572  (.I0(\edb_top_inst/n1762 ), .I1(\edb_top_inst/n1768 ), 
            .I2(\edb_top_inst/n1771 ), .I3(\edb_top_inst/n1780 ), .O(\edb_top_inst/n1781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3572 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3573  (.I0(\edb_top_inst/n1723 ), .I1(\edb_top_inst/n1741 ), 
            .I2(\edb_top_inst/n1758 ), .I3(\edb_top_inst/n1781 ), .O(\edb_top_inst/n1782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3573 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3574  (.I0(\edb_top_inst/la0/skip_count [14]), 
            .I1(\edb_top_inst/la0/skip_count [15]), .O(\edb_top_inst/n1783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3574 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3575  (.I0(\edb_top_inst/la0/skip_count [16]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16]), 
            .O(\edb_top_inst/n1784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3575 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3576  (.I0(\edb_top_inst/la0/skip_count [14]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14]), 
            .O(\edb_top_inst/n1785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3576 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3577  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/n1720 ), .O(\edb_top_inst/n1786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3577 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3578  (.I0(\edb_top_inst/n1783 ), .I1(\edb_top_inst/n1785 ), 
            .I2(\edb_top_inst/n1784 ), .I3(\edb_top_inst/n1786 ), .O(\edb_top_inst/n1787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3578 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3579  (.I0(\edb_top_inst/la0/skip_count [34]), 
            .I1(\edb_top_inst/n1767 ), .I2(\edb_top_inst/la0/skip_count [35]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35]), 
            .O(\edb_top_inst/n1788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb44b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3579 .LUTMASK = 16'hb44b;
    EFX_LUT4 \edb_top_inst/LUT__3580  (.I0(\edb_top_inst/n1733 ), .I1(\edb_top_inst/n1737 ), 
            .O(\edb_top_inst/n1789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3580 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3581  (.I0(\edb_top_inst/la0/skip_count [48]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48]), 
            .O(\edb_top_inst/n1790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3581 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3582  (.I0(\edb_top_inst/la0/skip_count [47]), 
            .I1(\edb_top_inst/n1732 ), .I2(\edb_top_inst/n1789 ), .I3(\edb_top_inst/n1790 ), 
            .O(\edb_top_inst/n1791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3582 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3583  (.I0(\edb_top_inst/n1787 ), .I1(\edb_top_inst/n1788 ), 
            .I2(\edb_top_inst/n1791 ), .O(\edb_top_inst/n1792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3583 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3584  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/la0/skip_count [56]), .I2(\edb_top_inst/la0/skip_count [57]), 
            .O(\edb_top_inst/n1793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3584 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3585  (.I0(\edb_top_inst/la0/skip_count [53]), 
            .I1(\edb_top_inst/la0/skip_count [54]), .I2(\edb_top_inst/n1743 ), 
            .I3(\edb_top_inst/n1793 ), .O(\edb_top_inst/n1794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3585 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3586  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/la0/skip_count [59]), .I2(\edb_top_inst/n1794 ), 
            .O(\edb_top_inst/n1795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3586 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3587  (.I0(\edb_top_inst/la0/skip_count [30]), 
            .I1(\edb_top_inst/n1746 ), .O(\edb_top_inst/n1796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3587 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3588  (.I0(\edb_top_inst/la0/skip_count [31]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31]), 
            .O(\edb_top_inst/n1797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3588 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3589  (.I0(\edb_top_inst/la0/skip_count [23]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .O(\edb_top_inst/n1798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3589 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3590  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/n1720 ), .I2(\edb_top_inst/n1725 ), .O(\edb_top_inst/n1799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3590 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3591  (.I0(\edb_top_inst/n1796 ), .I1(\edb_top_inst/n1798 ), 
            .I2(\edb_top_inst/n1797 ), .I3(\edb_top_inst/n1799 ), .O(\edb_top_inst/n1800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3591 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3592  (.I0(\edb_top_inst/la0/skip_count [60]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60]), 
            .O(\edb_top_inst/n1801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3592 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3593  (.I0(\edb_top_inst/n1739 ), .I1(\edb_top_inst/n1795 ), 
            .I2(\edb_top_inst/n1800 ), .I3(\edb_top_inst/n1801 ), .O(\edb_top_inst/n1802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3593 .LUTMASK = 16'h0708;
    EFX_LUT4 \edb_top_inst/LUT__3594  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/la0/skip_count [50]), .I2(\edb_top_inst/la0/skip_count [51]), 
            .O(\edb_top_inst/n1803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3594 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3595  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52]), 
            .I2(\edb_top_inst/n1803 ), .O(\edb_top_inst/n1804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3595 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__3596  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58]), 
            .I2(\edb_top_inst/n1794 ), .I3(\edb_top_inst/n1804 ), .O(\edb_top_inst/n1805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3596 .LUTMASK = 16'h6900;
    EFX_LUT4 \edb_top_inst/LUT__3597  (.I0(\edb_top_inst/la0/skip_count [52]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52]), 
            .I2(\edb_top_inst/la0/skip_count [58]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58]), 
            .O(\edb_top_inst/n1806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3597 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3598  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1738 ), 
            .I2(\edb_top_inst/n1803 ), .I3(\edb_top_inst/n1806 ), .O(\edb_top_inst/n1807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3598 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__3599  (.I0(\edb_top_inst/la0/skip_count [43]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43]), 
            .O(\edb_top_inst/n1808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3599 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3600  (.I0(\edb_top_inst/la0/skip_count [42]), 
            .I1(\edb_top_inst/n1732 ), .I2(\edb_top_inst/n1735 ), .I3(\edb_top_inst/n1808 ), 
            .O(\edb_top_inst/n1809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3600 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3601  (.I0(\edb_top_inst/n1739 ), .I1(\edb_top_inst/n1805 ), 
            .I2(\edb_top_inst/n1807 ), .I3(\edb_top_inst/n1809 ), .O(\edb_top_inst/n1810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3601 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3602  (.I0(\edb_top_inst/la0/skip_count [55]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55]), 
            .O(\edb_top_inst/n1811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3602 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3603  (.I0(\edb_top_inst/la0/skip_count [53]), 
            .I1(\edb_top_inst/la0/skip_count [54]), .I2(\edb_top_inst/n1743 ), 
            .O(\edb_top_inst/n1812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3603 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3604  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1738 ), 
            .I2(\edb_top_inst/n1812 ), .O(\edb_top_inst/n1813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3604 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3605  (.I0(\edb_top_inst/la0/skip_count [50]), 
            .I1(\edb_top_inst/la0/skip_count [51]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50]), 
            .O(\edb_top_inst/n1814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3605 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3606  (.I0(\edb_top_inst/la0/skip_count [50]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50]), 
            .I2(\edb_top_inst/la0/skip_count [51]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .O(\edb_top_inst/n1815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3606 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3607  (.I0(\edb_top_inst/la0/skip_count [49]), 
            .I1(\edb_top_inst/n1738 ), .O(\edb_top_inst/n1816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3607 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3608  (.I0(\edb_top_inst/n1814 ), .I1(\edb_top_inst/n1815 ), 
            .I2(\edb_top_inst/n1732 ), .I3(\edb_top_inst/n1816 ), .O(\edb_top_inst/n1817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3608 .LUTMASK = 16'ha333;
    EFX_LUT4 \edb_top_inst/LUT__3609  (.I0(\edb_top_inst/la0/skip_count [56]), 
            .I1(\edb_top_inst/la0/skip_count [57]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .O(\edb_top_inst/n1818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3609 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3610  (.I0(\edb_top_inst/la0/skip_count [56]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .I2(\edb_top_inst/la0/skip_count [57]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57]), 
            .O(\edb_top_inst/n1819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3610 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3611  (.I0(\edb_top_inst/n1818 ), .I1(\edb_top_inst/n1819 ), 
            .I2(\edb_top_inst/la0/skip_count [55]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55]), 
            .O(\edb_top_inst/n1820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a33, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3611 .LUTMASK = 16'h3a33;
    EFX_LUT4 \edb_top_inst/LUT__3612  (.I0(\edb_top_inst/n1817 ), .I1(\edb_top_inst/n1820 ), 
            .I2(\edb_top_inst/n1811 ), .I3(\edb_top_inst/n1813 ), .O(\edb_top_inst/n1821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3612 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__3613  (.I0(\edb_top_inst/n1792 ), .I1(\edb_top_inst/n1802 ), 
            .I2(\edb_top_inst/n1810 ), .I3(\edb_top_inst/n1821 ), .O(\edb_top_inst/n1822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3613 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3614  (.I0(\edb_top_inst/n1739 ), .I1(\edb_top_inst/n1743 ), 
            .I2(\edb_top_inst/la0/skip_count [53]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53]), 
            .O(\edb_top_inst/n1823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3614 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3615  (.I0(\edb_top_inst/n1751 ), .I1(\edb_top_inst/n1728 ), 
            .I2(\edb_top_inst/la0/skip_count [32]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32]), 
            .O(\edb_top_inst/n1824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3615 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3616  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1789 ), 
            .I2(\edb_top_inst/la0/skip_count [47]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47]), 
            .O(\edb_top_inst/n1825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3616 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3617  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/la0/skip_count [18]), .I2(\edb_top_inst/la0/skip_count [19]), 
            .I3(\edb_top_inst/n1721 ), .O(\edb_top_inst/n1826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3617 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3618  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1826 ), 
            .I2(\edb_top_inst/la0/skip_count [20]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20]), 
            .O(\edb_top_inst/n1827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3618 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3619  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1721 ), 
            .I2(\edb_top_inst/la0/skip_count [17]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17]), 
            .O(\edb_top_inst/n1828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3619 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3620  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/la0/skip_count [14]), .I2(\edb_top_inst/n1720 ), 
            .O(\edb_top_inst/n1829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3620 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3621  (.I0(\edb_top_inst/la0/skip_count [15]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15]), 
            .O(\edb_top_inst/n1830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3621 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3622  (.I0(\edb_top_inst/n1829 ), .I1(\edb_top_inst/n1830 ), 
            .I2(\edb_top_inst/n1827 ), .I3(\edb_top_inst/n1828 ), .O(\edb_top_inst/n1831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3622 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__3623  (.I0(\edb_top_inst/la0/skip_count [3]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3]), 
            .O(\edb_top_inst/n1832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3623 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3624  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .O(\edb_top_inst/n1833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3624 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3625  (.I0(\edb_top_inst/la0/skip_count [2]), 
            .I1(\edb_top_inst/n1832 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2]), 
            .I3(\edb_top_inst/n1833 ), .O(\edb_top_inst/n1834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3625 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3626  (.I0(\edb_top_inst/la0/skip_count [4]), 
            .I1(\edb_top_inst/n1717 ), .O(\edb_top_inst/n1835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3626 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3627  (.I0(\edb_top_inst/la0/skip_count [5]), 
            .I1(\edb_top_inst/n1835 ), .I2(\edb_top_inst/la0/skip_count [6]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6]), 
            .O(\edb_top_inst/n1836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb44b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3627 .LUTMASK = 16'hb44b;
    EFX_LUT4 \edb_top_inst/LUT__3628  (.I0(\edb_top_inst/la0/skip_count [13]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13]), 
            .I2(\edb_top_inst/n1720 ), .O(\edb_top_inst/n1837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3628 .LUTMASK = 16'h6969;
    EFX_LUT4 \edb_top_inst/LUT__3629  (.I0(\edb_top_inst/la0/skip_count [0]), 
            .I1(\edb_top_inst/la0/skip_count [1]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .O(\edb_top_inst/n1838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3629 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3630  (.I0(\edb_top_inst/n1838 ), .I1(\edb_top_inst/la0/skip_count [4]), 
            .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4]), 
            .I3(\edb_top_inst/n1717 ), .O(\edb_top_inst/n1839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3630 .LUTMASK = 16'h1441;
    EFX_LUT4 \edb_top_inst/LUT__3631  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8]), 
            .I2(\edb_top_inst/n1760 ), .I3(\edb_top_inst/n1839 ), .O(\edb_top_inst/n1840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3631 .LUTMASK = 16'h6900;
    EFX_LUT4 \edb_top_inst/LUT__3632  (.I0(\edb_top_inst/n1834 ), .I1(\edb_top_inst/n1836 ), 
            .I2(\edb_top_inst/n1837 ), .I3(\edb_top_inst/n1840 ), .O(\edb_top_inst/n1841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3632 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3633  (.I0(\edb_top_inst/la0/skip_count [5]), 
            .I1(\edb_top_inst/la0/skip_count [6]), .O(\edb_top_inst/n1842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3633 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3634  (.I0(\edb_top_inst/la0/skip_count [7]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7]), 
            .O(\edb_top_inst/n1843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3634 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3635  (.I0(\edb_top_inst/la0/skip_count [5]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5]), 
            .O(\edb_top_inst/n1844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3635 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3636  (.I0(\edb_top_inst/n1842 ), .I1(\edb_top_inst/n1844 ), 
            .I2(\edb_top_inst/n1843 ), .I3(\edb_top_inst/n1835 ), .O(\edb_top_inst/n1845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3636 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3637  (.I0(\edb_top_inst/la0/skip_count [17]), 
            .I1(\edb_top_inst/la0/skip_count [18]), .I2(\edb_top_inst/n1721 ), 
            .O(\edb_top_inst/n1846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3637 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3638  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1846 ), 
            .I2(\edb_top_inst/la0/skip_count [19]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19]), 
            .O(\edb_top_inst/n1847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3638 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3639  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22]), 
            .O(\edb_top_inst/n1848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3639 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3640  (.I0(\edb_top_inst/n1845 ), .I1(\edb_top_inst/n1848 ), 
            .I2(\edb_top_inst/n1751 ), .I3(\edb_top_inst/n1847 ), .O(\edb_top_inst/n1849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3640 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__3641  (.I0(\edb_top_inst/n1825 ), .I1(\edb_top_inst/n1831 ), 
            .I2(\edb_top_inst/n1841 ), .I3(\edb_top_inst/n1849 ), .O(\edb_top_inst/n1850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3641 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3642  (.I0(\edb_top_inst/la0/skip_count [22]), 
            .I1(\edb_top_inst/la0/skip_count [23]), .O(\edb_top_inst/n1851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3642 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3643  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1725 ), 
            .I2(\edb_top_inst/n1851 ), .O(\edb_top_inst/n1852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3643 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3644  (.I0(\edb_top_inst/la0/skip_count [25]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25]), 
            .O(\edb_top_inst/n1853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3644 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3645  (.I0(\edb_top_inst/la0/skip_count [24]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24]), 
            .I2(\edb_top_inst/n1852 ), .I3(\edb_top_inst/n1853 ), .O(\edb_top_inst/n1854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd6bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3645 .LUTMASK = 16'hd6bf;
    EFX_LUT4 \edb_top_inst/LUT__3646  (.I0(\edb_top_inst/la0/skip_count [38]), 
            .I1(\edb_top_inst/la0/skip_count [39]), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39]), 
            .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .O(\edb_top_inst/n1855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3646 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3647  (.I0(\edb_top_inst/la0/skip_count [38]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .I2(\edb_top_inst/la0/skip_count [39]), .I3(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39]), 
            .O(\edb_top_inst/n1856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3647 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3648  (.I0(\edb_top_inst/n1855 ), .I1(\edb_top_inst/n1856 ), 
            .I2(\edb_top_inst/n1730 ), .I3(\edb_top_inst/n1767 ), .O(\edb_top_inst/n1857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3648 .LUTMASK = 16'ha333;
    EFX_LUT4 \edb_top_inst/LUT__3649  (.I0(\edb_top_inst/la0/skip_count [12]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12]), 
            .O(\edb_top_inst/n1858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3649 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3650  (.I0(\edb_top_inst/la0/skip_count [8]), 
            .I1(\edb_top_inst/la0/skip_count [9]), .I2(\edb_top_inst/la0/skip_count [10]), 
            .I3(\edb_top_inst/n1760 ), .O(\edb_top_inst/n1859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3650 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3651  (.I0(\edb_top_inst/la0/skip_count [11]), 
            .I1(\edb_top_inst/n1858 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11]), 
            .I3(\edb_top_inst/n1859 ), .O(\edb_top_inst/n1860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3651 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3652  (.I0(\edb_top_inst/la0/skip_count [21]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21]), 
            .O(\edb_top_inst/n1861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3652 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3653  (.I0(\edb_top_inst/n1720 ), .I1(\edb_top_inst/n1721 ), 
            .I2(\edb_top_inst/n1724 ), .I3(\edb_top_inst/n1861 ), .O(\edb_top_inst/n1862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3653 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__3654  (.I0(\edb_top_inst/n1854 ), .I1(\edb_top_inst/n1857 ), 
            .I2(\edb_top_inst/n1860 ), .I3(\edb_top_inst/n1862 ), .O(\edb_top_inst/n1863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3654 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3655  (.I0(\edb_top_inst/n1823 ), .I1(\edb_top_inst/n1824 ), 
            .I2(\edb_top_inst/n1850 ), .I3(\edb_top_inst/n1863 ), .O(\edb_top_inst/n1864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3655 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3656  (.I0(\edb_top_inst/la0/skip_count [63]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63]), 
            .O(\edb_top_inst/n1865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3656 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3657  (.I0(\edb_top_inst/la0/skip_count [60]), 
            .I1(\edb_top_inst/la0/skip_count [61]), .O(\edb_top_inst/n1866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3657 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3658  (.I0(\edb_top_inst/n1732 ), .I1(\edb_top_inst/n1738 ), 
            .I2(\edb_top_inst/n1795 ), .I3(\edb_top_inst/n1866 ), .O(\edb_top_inst/n1867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3658 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3659  (.I0(\edb_top_inst/la0/skip_count [62]), 
            .I1(\edb_top_inst/n1865 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62]), 
            .I3(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3659 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3660  (.I0(\edb_top_inst/la0/skip_count [46]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .O(\edb_top_inst/n1869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3660 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3661  (.I0(\edb_top_inst/la0/skip_count [44]), 
            .I1(\edb_top_inst/n1732 ), .I2(\edb_top_inst/n1733 ), .O(\edb_top_inst/n1870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3661 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3662  (.I0(\edb_top_inst/la0/skip_count [45]), 
            .I1(\edb_top_inst/n1869 ), .I2(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45]), 
            .I3(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3662 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3663  (.I0(\edb_top_inst/la0/skip_count [59]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59]), 
            .O(\edb_top_inst/n1872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3663 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3664  (.I0(\edb_top_inst/la0/skip_count [58]), 
            .I1(\edb_top_inst/n1739 ), .I2(\edb_top_inst/n1794 ), .I3(\edb_top_inst/n1872 ), 
            .O(\edb_top_inst/n1873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3664 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3665  (.I0(\edb_top_inst/la0/skip_count [61]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61]), 
            .O(\edb_top_inst/n1874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3665 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3666  (.I0(\edb_top_inst/la0/skip_count [60]), 
            .I1(\edb_top_inst/n1739 ), .I2(\edb_top_inst/n1795 ), .I3(\edb_top_inst/n1874 ), 
            .O(\edb_top_inst/n1875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3666 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3667  (.I0(\edb_top_inst/n1868 ), .I1(\edb_top_inst/n1871 ), 
            .I2(\edb_top_inst/n1873 ), .I3(\edb_top_inst/n1875 ), .O(\edb_top_inst/n1876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3667 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3668  (.I0(\edb_top_inst/n1782 ), .I1(\edb_top_inst/n1822 ), 
            .I2(\edb_top_inst/n1864 ), .I3(\edb_top_inst/n1876 ), .O(\edb_top_inst/n1877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3668 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3669  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .I1(\edb_top_inst/n1877 ), .O(\edb_top_inst/la0/trigger_skipper_n/n138 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3669 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3670  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/n1877 ), .O(\edb_top_inst/la0/trigger_skipper_n/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3670 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3671  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [1]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3671 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3672  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [2]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3672 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3673  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [3]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3673 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3674  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [4]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3674 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3675  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [5]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3675 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3676  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [6]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3676 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3677  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [7]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3677 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3678  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [8]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3678 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3679  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [9]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3679 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3680  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [10]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3680 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3681  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [11]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3681 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3682  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [12]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3682 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3683  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [13]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3683 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3684  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [14]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3684 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3685  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [15]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3685 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3686  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [16]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3686 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3687  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [17]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3687 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3688  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [18]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3688 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3689  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [19]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3689 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3690  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [20]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3690 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3691  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [21]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3691 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3692  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [22]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3692 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3693  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [23]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3693 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3694  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [24]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3694 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3695  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [25]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3695 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3696  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [26]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3696 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3697  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [27]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3697 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3698  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [28]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3698 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3699  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [29]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3699 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3700  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [30]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3700 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3701  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [31]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3701 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3702  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [32]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3702 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3703  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [33]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3703 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3704  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [34]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3704 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3705  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [35]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3705 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3706  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [36]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3706 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3707  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [37]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3707 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3708  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [38]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3708 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3709  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [39]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3709 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3710  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [40]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3710 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3711  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [41]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3711 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3712  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [42]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3712 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3713  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [43]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3713 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3714  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [44]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3714 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3715  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [45]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3715 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3716  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [46]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3716 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3717  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [47]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3717 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3718  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [48]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3718 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3719  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [49]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3719 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3720  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [50]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3720 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3721  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [51]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3721 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3722  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [52]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3722 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3723  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [53]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3723 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3724  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [54]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3724 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3725  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [55]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3725 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3726  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [56]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3726 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3727  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [57]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3727 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3728  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [58]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3728 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3729  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [59]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3729 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3730  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [60]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3730 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3731  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [61]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3731 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3732  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [62]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3732 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3733  (.I0(\edb_top_inst/n1877 ), .I1(\edb_top_inst/la0/trigger_skipper_n/n73 [63]), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n138 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3733 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3734  (.I0(\edb_top_inst/la0/ts_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n1878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3734 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3735  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n1879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3735 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3736  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n1880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3736 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3737  (.I0(\edb_top_inst/n1880 ), .I1(\edb_top_inst/n1879 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [5]), .I3(\edb_top_inst/la0/la_trig_pos [1]), 
            .O(\edb_top_inst/n1881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hebd5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3737 .LUTMASK = 16'hebd5;
    EFX_LUT4 \edb_top_inst/LUT__3738  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n1882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3738 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3739  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n1883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3739 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3740  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1882 ), .I2(\edb_top_inst/n1883 ), .I3(\edb_top_inst/la0/la_trig_pos [6]), 
            .O(\edb_top_inst/n1884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h708f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3740 .LUTMASK = 16'h708f;
    EFX_LUT4 \edb_top_inst/LUT__3741  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [7]), .I2(\edb_top_inst/la0/la_trig_pos [3]), 
            .I3(\edb_top_inst/n1883 ), .O(\edb_top_inst/n1885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3741 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3742  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n1886 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3742 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3743  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1886 ), .I2(\edb_top_inst/n1883 ), .I3(\edb_top_inst/la0/la_trig_pos [4]), 
            .O(\edb_top_inst/n1887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd02f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3743 .LUTMASK = 16'hd02f;
    EFX_LUT4 \edb_top_inst/LUT__3744  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n1888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3744 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3745  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/n1888 ), .O(\edb_top_inst/n1889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3745 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3746  (.I0(\edb_top_inst/n1889 ), .I1(\edb_top_inst/la0/la_trig_pos [15]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/la0/la_trig_pos [13]), 
            .O(\edb_top_inst/n1890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3746 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__3747  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .O(\edb_top_inst/n1891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3747 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3748  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/n1891 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n1892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3748 .LUTMASK = 16'hf20d;
    EFX_LUT4 \edb_top_inst/LUT__3749  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .O(\edb_top_inst/n1893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3749 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3750  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/n1893 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [2]), .O(\edb_top_inst/n1894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3750 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3751  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n1895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3751 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3752  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [0]), .I2(\edb_top_inst/n1895 ), 
            .I3(\edb_top_inst/la0/la_trig_pos [16]), .O(\edb_top_inst/n1896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f8a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3752 .LUTMASK = 16'h7f8a;
    EFX_LUT4 \edb_top_inst/LUT__3753  (.I0(\edb_top_inst/n1886 ), .I1(\edb_top_inst/n1893 ), 
            .I2(\edb_top_inst/n1896 ), .I3(\edb_top_inst/la0/la_trig_pos [0]), 
            .O(\edb_top_inst/n1897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3753 .LUTMASK = 16'h0708;
    EFX_LUT4 \edb_top_inst/LUT__3754  (.I0(\edb_top_inst/n1890 ), .I1(\edb_top_inst/n1894 ), 
            .I2(\edb_top_inst/n1892 ), .I3(\edb_top_inst/n1897 ), .O(\edb_top_inst/n1898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3754 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3755  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .O(\edb_top_inst/n1899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3755 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3756  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/n1899 ), .O(\edb_top_inst/n1900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3756 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3757  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/n1888 ), .O(\edb_top_inst/n1901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3757 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3758  (.I0(\edb_top_inst/n1900 ), .I1(\edb_top_inst/n1901 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [12]), .I3(\edb_top_inst/la0/la_trig_pos [11]), 
            .O(\edb_top_inst/n1902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3758 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__3759  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n1903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3759 .LUTMASK = 16'hfe00;
    EFX_LUT4 \edb_top_inst/LUT__3760  (.I0(\edb_top_inst/n1888 ), .I1(\edb_top_inst/n1882 ), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n1904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3760 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3761  (.I0(\edb_top_inst/n1903 ), .I1(\edb_top_inst/la0/la_trig_pos [14]), 
            .I2(\edb_top_inst/la0/la_trig_pos [8]), .I3(\edb_top_inst/n1904 ), 
            .O(\edb_top_inst/n1905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3761 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3762  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1882 ), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .I3(\edb_top_inst/la0/la_window_depth [4]), .O(\edb_top_inst/n1906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3762 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__3763  (.I0(\edb_top_inst/n1902 ), .I1(\edb_top_inst/n1905 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [10]), .I3(\edb_top_inst/n1906 ), 
            .O(\edb_top_inst/n1907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3763 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__3764  (.I0(\edb_top_inst/n1885 ), .I1(\edb_top_inst/n1887 ), 
            .I2(\edb_top_inst/n1898 ), .I3(\edb_top_inst/n1907 ), .O(\edb_top_inst/n1908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3764 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3765  (.I0(\edb_top_inst/n1881 ), .I1(\edb_top_inst/n1884 ), 
            .I2(\edb_top_inst/n1908 ), .O(\edb_top_inst/n1909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3765 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3766  (.I0(\edb_top_inst/n1878 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .O(\edb_top_inst/n1910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3766 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__3767  (.I0(\edb_top_inst/n1909 ), .I1(\edb_top_inst/n1878 ), 
            .I2(\edb_top_inst/n1910 ), .O(\edb_top_inst/n1911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3767 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__3768  (.I0(\edb_top_inst/la0/la_trig_pos [13]), 
            .I1(\edb_top_inst/la0/la_trig_pos [14]), .I2(\edb_top_inst/la0/la_trig_pos [15]), 
            .I3(\edb_top_inst/la0/la_trig_pos [16]), .O(\edb_top_inst/n1912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3768 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3769  (.I0(\edb_top_inst/la0/la_trig_pos [10]), 
            .I1(\edb_top_inst/la0/la_trig_pos [11]), .I2(\edb_top_inst/la0/la_trig_pos [12]), 
            .I3(\edb_top_inst/n1912 ), .O(\edb_top_inst/n1913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3769 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3770  (.I0(\edb_top_inst/la0/la_trig_pos [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [4]), .I2(\edb_top_inst/la0/la_trig_pos [5]), 
            .I3(\edb_top_inst/la0/la_trig_pos [6]), .O(\edb_top_inst/n1914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3770 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3771  (.I0(\edb_top_inst/la0/la_trig_pos [3]), 
            .I1(\edb_top_inst/la0/la_trig_pos [7]), .O(\edb_top_inst/n1915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3771 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3772  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_trig_pos [1]), .I2(\edb_top_inst/la0/la_trig_pos [8]), 
            .I3(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n1916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3772 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3773  (.I0(\edb_top_inst/n1913 ), .I1(\edb_top_inst/n1914 ), 
            .I2(\edb_top_inst/n1915 ), .I3(\edb_top_inst/n1916 ), .O(\edb_top_inst/n1917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3773 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3774  (.I0(\edb_top_inst/la0/la_num_trigger [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), .O(\edb_top_inst/n1918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3774 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3775  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .I2(\edb_top_inst/la0/la_num_trigger [2]), 
            .I3(\edb_top_inst/la0/la_num_trigger [3]), .O(\edb_top_inst/n1919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3775 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3776  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/la0/la_num_trigger [5]), .I2(\edb_top_inst/la0/la_num_trigger [6]), 
            .O(\edb_top_inst/n1920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3776 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3777  (.I0(\edb_top_inst/n1919 ), .I1(\edb_top_inst/n1920 ), 
            .O(\edb_top_inst/n1921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3777 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3778  (.I0(\edb_top_inst/la0/la_num_trigger [7]), 
            .I1(\edb_top_inst/n1918 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I3(\edb_top_inst/n1921 ), .O(\edb_top_inst/n1922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3778 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3779  (.I0(\edb_top_inst/la0/la_num_trigger [7]), 
            .I1(\edb_top_inst/la0/la_num_trigger [8]), .I2(\edb_top_inst/n1919 ), 
            .I3(\edb_top_inst/n1920 ), .O(\edb_top_inst/n1923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3779 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3780  (.I0(\edb_top_inst/la0/la_num_trigger [9]), 
            .I1(\edb_top_inst/la0/la_num_trigger [10]), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I3(\edb_top_inst/n1923 ), .O(\edb_top_inst/n1924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3780 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__3781  (.I0(\edb_top_inst/la0/la_num_trigger [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), .O(\edb_top_inst/n1925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3781 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3782  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/n1919 ), .O(\edb_top_inst/n1926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3782 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3783  (.I0(\edb_top_inst/la0/la_num_trigger [5]), 
            .I1(\edb_top_inst/n1925 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I3(\edb_top_inst/n1926 ), .O(\edb_top_inst/n1927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3783 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3784  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .O(\edb_top_inst/n1928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3784 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3785  (.I0(\edb_top_inst/la0/la_num_trigger [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), .O(\edb_top_inst/n1929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3785 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3786  (.I0(\edb_top_inst/la0/la_num_trigger [0]), 
            .I1(\edb_top_inst/la0/la_num_trigger [1]), .O(\edb_top_inst/n1930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3786 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3787  (.I0(\edb_top_inst/la0/la_num_trigger [2]), 
            .I1(\edb_top_inst/n1929 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I3(\edb_top_inst/n1930 ), .O(\edb_top_inst/n1931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3787 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3788  (.I0(\edb_top_inst/la0/la_num_trigger [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), .I2(\edb_top_inst/n1919 ), 
            .O(\edb_top_inst/n1932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3788 .LUTMASK = 16'h6969;
    EFX_LUT4 \edb_top_inst/LUT__3789  (.I0(\edb_top_inst/la0/la_num_trigger [11]), 
            .I1(\edb_top_inst/la0/la_num_trigger [13]), .I2(\edb_top_inst/la0/la_num_trigger [14]), 
            .I3(\edb_top_inst/la0/la_num_trigger [15]), .O(\edb_top_inst/n1933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3789 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3790  (.I0(\edb_top_inst/la0/la_num_trigger [12]), 
            .I1(\edb_top_inst/la0/la_num_trigger [16]), .I2(\edb_top_inst/n1933 ), 
            .O(\edb_top_inst/n1934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3790 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3791  (.I0(\edb_top_inst/n1928 ), .I1(\edb_top_inst/n1931 ), 
            .I2(\edb_top_inst/n1932 ), .I3(\edb_top_inst/n1934 ), .O(\edb_top_inst/n1935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3791 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3792  (.I0(\edb_top_inst/n1922 ), .I1(\edb_top_inst/n1924 ), 
            .I2(\edb_top_inst/n1927 ), .I3(\edb_top_inst/n1935 ), .O(\edb_top_inst/n1936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3792 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3793  (.I0(\edb_top_inst/n1917 ), .I1(\edb_top_inst/n1936 ), 
            .O(\edb_top_inst/n1937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3793 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3794  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_window_depth [4]), .I2(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n1938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3794 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3795  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/n1938 ), 
            .O(\edb_top_inst/n1939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3795 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3796  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [3]), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/n1891 ), .O(\edb_top_inst/n1940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3796 .LUTMASK = 16'h0e03;
    EFX_LUT4 \edb_top_inst/LUT__3797  (.I0(\edb_top_inst/la0/la_trig_pos [9]), 
            .I1(\edb_top_inst/la0/la_trig_pos [10]), .I2(\edb_top_inst/n1939 ), 
            .I3(\edb_top_inst/n1940 ), .O(\edb_top_inst/n1941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3797 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__3798  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/n1888 ), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .I3(\edb_top_inst/la0/la_trig_pos [14]), .O(\edb_top_inst/n1942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4cbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3798 .LUTMASK = 16'h4cbf;
    EFX_LUT4 \edb_top_inst/LUT__3799  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_trig_pos [14]), 
            .I3(\edb_top_inst/n1888 ), .O(\edb_top_inst/n1943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3799 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3800  (.I0(\edb_top_inst/n1901 ), .I1(\edb_top_inst/n1942 ), 
            .I2(\edb_top_inst/n1943 ), .I3(\edb_top_inst/la0/la_trig_pos [13]), 
            .O(\edb_top_inst/n1944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3800 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__3801  (.I0(\edb_top_inst/n1886 ), .I1(\edb_top_inst/n1888 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [12]), .O(\edb_top_inst/n1945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3801 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3802  (.I0(\edb_top_inst/n1895 ), .I1(\edb_top_inst/n1945 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [15]), .I3(\edb_top_inst/la0/la_window_depth [4]), 
            .O(\edb_top_inst/n1946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdff3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3802 .LUTMASK = 16'hdff3;
    EFX_LUT4 \edb_top_inst/LUT__3803  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_window_depth [1]), .I2(\edb_top_inst/la0/la_window_depth [2]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n1947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3803 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3804  (.I0(\edb_top_inst/la0/la_trig_pos [16]), 
            .I1(\edb_top_inst/n1947 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .O(\edb_top_inst/n1948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9e9e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3804 .LUTMASK = 16'h9e9e;
    EFX_LUT4 \edb_top_inst/LUT__3805  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_trig_pos [3]), .I2(\edb_top_inst/n1893 ), 
            .O(\edb_top_inst/n1949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3805 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__3806  (.I0(\edb_top_inst/n1948 ), .I1(\edb_top_inst/la0/la_trig_pos [11]), 
            .I2(\edb_top_inst/n1901 ), .I3(\edb_top_inst/n1949 ), .O(\edb_top_inst/n1950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3806 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__3807  (.I0(\edb_top_inst/n1941 ), .I1(\edb_top_inst/n1944 ), 
            .I2(\edb_top_inst/n1946 ), .I3(\edb_top_inst/n1950 ), .O(\edb_top_inst/n1951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3807 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3808  (.I0(\edb_top_inst/n1886 ), .I1(\edb_top_inst/n1938 ), 
            .O(\edb_top_inst/n1952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3808 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3809  (.I0(\edb_top_inst/n1891 ), .I1(\edb_top_inst/la0/la_window_depth [0]), 
            .I2(\edb_top_inst/n1883 ), .O(\edb_top_inst/n1953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3809 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__3810  (.I0(\edb_top_inst/n1952 ), .I1(\edb_top_inst/n1953 ), 
            .I2(\edb_top_inst/la0/la_trig_pos [8]), .I3(\edb_top_inst/la0/la_trig_pos [7]), 
            .O(\edb_top_inst/n1954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3810 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__3811  (.I0(\edb_top_inst/n1894 ), .I1(\edb_top_inst/n1887 ), 
            .O(\edb_top_inst/n1955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3811 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3812  (.I0(\edb_top_inst/n1954 ), .I1(\edb_top_inst/n1884 ), 
            .I2(\edb_top_inst/n1881 ), .I3(\edb_top_inst/n1955 ), .O(\edb_top_inst/n1956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3812 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3813  (.I0(\edb_top_inst/n1903 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), .I3(\edb_top_inst/n1906 ), 
            .O(\edb_top_inst/n1957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3813 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3814  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/n1891 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), .O(\edb_top_inst/n1958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3814 .LUTMASK = 16'hf20d;
    EFX_LUT4 \edb_top_inst/LUT__3815  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1882 ), .I2(\edb_top_inst/n1883 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .O(\edb_top_inst/n1959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h708f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3815 .LUTMASK = 16'h708f;
    EFX_LUT4 \edb_top_inst/LUT__3816  (.I0(\edb_top_inst/n1886 ), .I1(\edb_top_inst/n1893 ), 
            .I2(\edb_top_inst/n1959 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
            .O(\edb_top_inst/n1960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3816 .LUTMASK = 16'h0708;
    EFX_LUT4 \edb_top_inst/LUT__3817  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/n1883 ), .O(\edb_top_inst/n1961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3817 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3818  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/n1893 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), .O(\edb_top_inst/n1962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3818 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3819  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1886 ), .I2(\edb_top_inst/n1883 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .O(\edb_top_inst/n1963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd02f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3819 .LUTMASK = 16'hd02f;
    EFX_LUT4 \edb_top_inst/LUT__3820  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), .I2(\edb_top_inst/n1879 ), 
            .I3(\edb_top_inst/n1880 ), .O(\edb_top_inst/n1964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3820 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__3821  (.I0(\edb_top_inst/n1961 ), .I1(\edb_top_inst/n1962 ), 
            .I2(\edb_top_inst/n1963 ), .I3(\edb_top_inst/n1964 ), .O(\edb_top_inst/n1965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3821 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3822  (.I0(\edb_top_inst/n1957 ), .I1(\edb_top_inst/n1958 ), 
            .I2(\edb_top_inst/n1960 ), .I3(\edb_top_inst/n1965 ), .O(\edb_top_inst/n1966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3822 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3823  (.I0(\edb_top_inst/n1886 ), .I1(\edb_top_inst/n1882 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n1883 ), 
            .O(\edb_top_inst/n1967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3823 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3824  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/n1967 ), .O(\edb_top_inst/n1968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3824 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3825  (.I0(\edb_top_inst/la0/la_window_depth [2]), 
            .I1(\edb_top_inst/n1882 ), .I2(\edb_top_inst/la0/la_window_depth [4]), 
            .I3(\edb_top_inst/la0/la_window_depth [3]), .O(\edb_top_inst/n1969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h010e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3825 .LUTMASK = 16'h010e;
    EFX_LUT4 \edb_top_inst/LUT__3826  (.I0(\edb_top_inst/n1969 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), .I3(\edb_top_inst/n1953 ), 
            .O(\edb_top_inst/n1970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3826 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3827  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/n1939 ), .I3(\edb_top_inst/n1940 ), .O(\edb_top_inst/n1971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3827 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__3828  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), .O(\edb_top_inst/n1972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3828 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3829  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/n1891 ), .I2(\edb_top_inst/n1879 ), .I3(\edb_top_inst/n1972 ), 
            .O(\edb_top_inst/n1973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3829 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__3830  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_window_depth [0]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I3(\edb_top_inst/la0/la_window_depth [2]), .O(\edb_top_inst/n1974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbef1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3830 .LUTMASK = 16'hbef1;
    EFX_LUT4 \edb_top_inst/LUT__3831  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), 
            .I1(\edb_top_inst/n1974 ), .I2(\edb_top_inst/n1883 ), .O(\edb_top_inst/n1975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3831 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3832  (.I0(\edb_top_inst/la0/la_window_depth [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I3(\edb_top_inst/n1880 ), .O(\edb_top_inst/n1976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdcf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3832 .LUTMASK = 16'hbdcf;
    EFX_LUT4 \edb_top_inst/LUT__3833  (.I0(\edb_top_inst/la0/la_window_depth [4]), 
            .I1(\edb_top_inst/n1903 ), .I2(\edb_top_inst/n1947 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .O(\edb_top_inst/n1977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3833 .LUTMASK = 16'hfe01;
    EFX_LUT4 \edb_top_inst/LUT__3834  (.I0(\edb_top_inst/n1975 ), .I1(\edb_top_inst/n1973 ), 
            .I2(\edb_top_inst/n1976 ), .I3(\edb_top_inst/n1977 ), .O(\edb_top_inst/n1978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3834 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__3835  (.I0(\edb_top_inst/n1968 ), .I1(\edb_top_inst/n1970 ), 
            .I2(\edb_top_inst/n1971 ), .I3(\edb_top_inst/n1978 ), .O(\edb_top_inst/n1979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3835 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3836  (.I0(\edb_top_inst/n1956 ), .I1(\edb_top_inst/n1966 ), 
            .I2(\edb_top_inst/n1951 ), .I3(\edb_top_inst/n1979 ), .O(\edb_top_inst/n1980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3836 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__3837  (.I0(\edb_top_inst/n1980 ), .I1(\edb_top_inst/n1937 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .O(\edb_top_inst/n1981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3837 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__3838  (.I0(\edb_top_inst/n1936 ), .I1(\edb_top_inst/n1878 ), 
            .I2(\edb_top_inst/n1966 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .O(\edb_top_inst/n1982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3838 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__3839  (.I0(\edb_top_inst/n1981 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I2(\edb_top_inst/n1982 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n1983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3839 .LUTMASK = 16'hf0bb;
    EFX_LUT4 \edb_top_inst/LUT__3840  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), 
            .I1(\edb_top_inst/la0/la_trig_pos [2]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I3(\edb_top_inst/la0/la_trig_pos [3]), .O(\edb_top_inst/n1984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3840 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3841  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), 
            .I1(\edb_top_inst/la0/la_trig_pos [5]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I3(\edb_top_inst/la0/la_trig_pos [9]), .O(\edb_top_inst/n1985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3841 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3842  (.I0(\edb_top_inst/la0/la_trig_pos [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I3(\edb_top_inst/la0/la_trig_pos [1]), .O(\edb_top_inst/n1986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3842 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3843  (.I0(\edb_top_inst/n1913 ), .I1(\edb_top_inst/n1984 ), 
            .I2(\edb_top_inst/n1985 ), .I3(\edb_top_inst/n1986 ), .O(\edb_top_inst/n1987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3843 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3844  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I1(\edb_top_inst/la0/la_trig_pos [4]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I3(\edb_top_inst/la0/la_trig_pos [7]), .O(\edb_top_inst/n1988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3844 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3845  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .I1(\edb_top_inst/la0/la_trig_pos [6]), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .I3(\edb_top_inst/la0/la_trig_pos [8]), .O(\edb_top_inst/n1989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3845 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3846  (.I0(\edb_top_inst/n1987 ), .I1(\edb_top_inst/n1988 ), 
            .I2(\edb_top_inst/n1989 ), .O(\edb_top_inst/n1990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3846 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3847  (.I0(\edb_top_inst/n1990 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .O(\edb_top_inst/n1991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3847 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3848  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I3(\edb_top_inst/n1917 ), .O(\edb_top_inst/n1992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3848 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__3849  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n1993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3849 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3850  (.I0(\edb_top_inst/n1992 ), .I1(\edb_top_inst/n1991 ), 
            .I2(\edb_top_inst/n1993 ), .O(\edb_top_inst/n1994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3850 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__3851  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .O(\edb_top_inst/n1995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3851 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3852  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n1996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3852 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3853  (.I0(\edb_top_inst/n1966 ), .I1(\edb_top_inst/n1878 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .I3(\edb_top_inst/n1996 ), 
            .O(\edb_top_inst/n1997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3853 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3854  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/n1990 ), .I2(\edb_top_inst/n1995 ), .I3(\edb_top_inst/n1997 ), 
            .O(\edb_top_inst/n1998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3854 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__3855  (.I0(\edb_top_inst/n1983 ), .I1(\edb_top_inst/n1911 ), 
            .I2(\edb_top_inst/n1994 ), .I3(\edb_top_inst/n1998 ), .O(\edb_top_inst/la0/la_biu_inst/next_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3855 .LUTMASK = 16'he0ff;
    EFX_LUT4 \edb_top_inst/LUT__3856  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), .O(\edb_top_inst/la0/la_biu_inst/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3856 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3857  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/n1481 ), .O(\edb_top_inst/la0/la_biu_inst/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3857 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3858  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), .O(\edb_top_inst/la0/la_biu_inst/n1248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3858 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3859  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3859 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__3860  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/n1832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3860 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3861  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .O(\edb_top_inst/n1999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3861 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3862  (.I0(\edb_top_inst/n1878 ), .I1(\edb_top_inst/n1999 ), 
            .I2(\edb_top_inst/n1909 ), .O(\edb_top_inst/n2000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3862 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3863  (.I0(\edb_top_inst/n2000 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/n1983 ), .O(\edb_top_inst/la0/la_biu_inst/n1214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3863 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__3864  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [3]), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n5970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3864 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3865  (.I0(\edb_top_inst/n1909 ), .I1(\edb_top_inst/n1936 ), 
            .I2(\edb_top_inst/la0/la_stop_trig ), .I3(\edb_top_inst/n1878 ), 
            .O(\edb_top_inst/n2001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3865 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__3866  (.I0(\edb_top_inst/n1878 ), .I1(\edb_top_inst/n1936 ), 
            .I2(\edb_top_inst/n1966 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .O(\edb_top_inst/n2002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3866 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__3867  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/n2002 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .O(\edb_top_inst/n2003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3867 .LUTMASK = 16'h8787;
    EFX_LUT4 \edb_top_inst/LUT__3868  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I2(\edb_top_inst/n2003 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), .O(\edb_top_inst/n2004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedfb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3868 .LUTMASK = 16'hedfb;
    EFX_LUT4 \edb_top_inst/LUT__3869  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I1(\edb_top_inst/n1993 ), .O(\edb_top_inst/n2005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3869 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3870  (.I0(\edb_top_inst/n1980 ), .I1(\edb_top_inst/n1937 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I3(\edb_top_inst/n2005 ), 
            .O(\edb_top_inst/n2006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3870 .LUTMASK = 16'heff0;
    EFX_LUT4 \edb_top_inst/LUT__3871  (.I0(\edb_top_inst/n2001 ), .I1(\edb_top_inst/n2004 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I3(\edb_top_inst/n2006 ), 
            .O(\edb_top_inst/la0/la_biu_inst/next_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h37f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3871 .LUTMASK = 16'h37f3;
    EFX_LUT4 \edb_top_inst/LUT__3872  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), .I2(\edb_top_inst/n1917 ), 
            .O(\edb_top_inst/n2007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3872 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__3873  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/n2007 ), .I2(\edb_top_inst/n1991 ), .I3(\edb_top_inst/n1993 ), 
            .O(\edb_top_inst/n2008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3873 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3874  (.I0(\edb_top_inst/n1936 ), .I1(\edb_top_inst/n1917 ), 
            .I2(\edb_top_inst/n1980 ), .O(\edb_top_inst/n2009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3874 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3875  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/n2009 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/n2008 ), .O(\edb_top_inst/n2010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3875 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3876  (.I0(\edb_top_inst/n1878 ), .I1(\edb_top_inst/n1909 ), 
            .I2(\edb_top_inst/n1936 ), .I3(\edb_top_inst/n1910 ), .O(\edb_top_inst/n2011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3876 .LUTMASK = 16'hbe00;
    EFX_LUT4 \edb_top_inst/LUT__3877  (.I0(\edb_top_inst/n1966 ), .I1(\edb_top_inst/n1878 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .O(\edb_top_inst/n2012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3877 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__3878  (.I0(\edb_top_inst/n1990 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .I3(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .O(\edb_top_inst/n2013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3878 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__3879  (.I0(\edb_top_inst/n2012 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I2(\edb_top_inst/n1993 ), .I3(\edb_top_inst/n2013 ), .O(\edb_top_inst/n2014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3879 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3880  (.I0(\edb_top_inst/n2011 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I2(\edb_top_inst/n2010 ), .I3(\edb_top_inst/n2014 ), .O(\edb_top_inst/la0/la_biu_inst/next_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3880 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3881  (.I0(\edb_top_inst/la0/la_biu_inst/n335 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
            .O(\edb_top_inst/ceg_net18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3881 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__3882  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3882 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3883  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [0]), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state [1]), 
            .O(\edb_top_inst/ceg_net24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3883 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3884  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .I2(\edb_top_inst/n1999 ), 
            .O(\edb_top_inst/n2015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3884 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3885  (.I0(\edb_top_inst/n1878 ), .I1(\edb_top_inst/n2015 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3885 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__3886  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [0]), .I2(\edb_top_inst/la0/la_biu_inst/curr_state [1]), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state [3]), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3886 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__3887  (.I0(\edb_top_inst/la0/la_biu_inst/n1839 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n2016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3887 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3888  (.I0(\edb_top_inst/n1966 ), .I1(\edb_top_inst/n2016 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3888 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3889  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state [1]), .I2(\edb_top_inst/n1993 ), 
            .I3(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3889 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__3890  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3890 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3891  (.I0(\edb_top_inst/n2016 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/~ceg_net27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3891 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3892  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n1547 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3892 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3893  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [0]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [15]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3893 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3894  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [16]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3894 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3895  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [17]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3895 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3896  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [18]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3896 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3897  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [19]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3897 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3898  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [5]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [20]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3898 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3899  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [21]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3899 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3900  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [7]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [22]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3900 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3901  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [23]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3901 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3902  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg [24]), .I2(\edb_top_inst/n1547 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3902 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3903  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), 
            .I1(\edb_top_inst/n1886 ), .O(\edb_top_inst/n2017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3903 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3904  (.I0(\edb_top_inst/n1893 ), .I1(\edb_top_inst/n2017 ), 
            .O(\edb_top_inst/n2018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3904 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3905  (.I0(\edb_top_inst/n1947 ), .I1(\edb_top_inst/n1906 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
            .I3(\edb_top_inst/n2018 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3905 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3906  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .I2(\edb_top_inst/la0/la_window_depth [0]), 
            .O(\edb_top_inst/n2019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3906 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3907  (.I0(\edb_top_inst/n2019 ), .I1(\edb_top_inst/n1880 ), 
            .O(\edb_top_inst/n2020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3907 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3908  (.I0(\edb_top_inst/n1895 ), .I1(\edb_top_inst/n1906 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1]), 
            .I3(\edb_top_inst/n2020 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3908 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3909  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3909 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3910  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), .I2(\edb_top_inst/n2021 ), 
            .I3(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3910 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3911  (.I0(\edb_top_inst/n2022 ), .I1(\edb_top_inst/n1893 ), 
            .O(\edb_top_inst/n2023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3911 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3912  (.I0(\edb_top_inst/n1969 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2]), 
            .I2(\edb_top_inst/n2023 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3912 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3913  (.I0(\edb_top_inst/la0/la_window_depth [3]), 
            .I1(\edb_top_inst/la0/la_window_depth [2]), .I2(\edb_top_inst/n1906 ), 
            .O(\edb_top_inst/n2024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3913 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__3914  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), .I2(\edb_top_inst/la0/la_window_depth [0]), 
            .O(\edb_top_inst/n2025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3914 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3915  (.I0(\edb_top_inst/n2025 ), .I1(\edb_top_inst/n2019 ), 
            .I2(\edb_top_inst/la0/la_window_depth [1]), .O(\edb_top_inst/n2026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3915 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3916  (.I0(\edb_top_inst/n2026 ), .I1(\edb_top_inst/n1893 ), 
            .O(\edb_top_inst/n2027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3916 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3917  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3]), 
            .I1(\edb_top_inst/n2024 ), .I2(\edb_top_inst/n2027 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3917 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3918  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3918 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3919  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3919 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3920  (.I0(\edb_top_inst/n2029 ), .I1(\edb_top_inst/n2028 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3920 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3921  (.I0(\edb_top_inst/n2030 ), .I1(\edb_top_inst/n2017 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n1883 ), 
            .O(\edb_top_inst/n2031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3921 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3922  (.I0(\edb_top_inst/n1900 ), .I1(\edb_top_inst/n2024 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4]), 
            .I3(\edb_top_inst/n2031 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3922 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3923  (.I0(\edb_top_inst/la0/la_window_depth [1]), 
            .I1(\edb_top_inst/n2019 ), .O(\edb_top_inst/n2032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3923 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3924  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3924 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3925  (.I0(\edb_top_inst/n2033 ), .I1(\edb_top_inst/n2029 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3925 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3926  (.I0(\edb_top_inst/n2034 ), .I1(\edb_top_inst/n2032 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n1883 ), 
            .O(\edb_top_inst/n2035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3926 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3927  (.I0(\edb_top_inst/n1899 ), .I1(\edb_top_inst/n2024 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5]), 
            .I3(\edb_top_inst/n2035 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3927 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3928  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/la0/la_window_depth [3]), 
            .I2(\edb_top_inst/n2024 ), .O(\edb_top_inst/n2036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3928 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__3929  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3929 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3930  (.I0(\edb_top_inst/n2037 ), .I1(\edb_top_inst/n2033 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3930 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3931  (.I0(\edb_top_inst/n2038 ), .I1(\edb_top_inst/n2022 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n1883 ), 
            .O(\edb_top_inst/n2039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3931 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3932  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6]), 
            .I1(\edb_top_inst/n2036 ), .I2(\edb_top_inst/n2039 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3932 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3933  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3933 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3934  (.I0(\edb_top_inst/n2040 ), .I1(\edb_top_inst/n2037 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3934 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3935  (.I0(\edb_top_inst/n2041 ), .I1(\edb_top_inst/n2026 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/n1883 ), 
            .O(\edb_top_inst/n2042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3935 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3936  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/n1938 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7]), 
            .I3(\edb_top_inst/n2042 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3936 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3937  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3937 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3938  (.I0(\edb_top_inst/n2043 ), .I1(\edb_top_inst/n2040 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3938 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3939  (.I0(\edb_top_inst/n2044 ), .I1(\edb_top_inst/n2017 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3939 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__3940  (.I0(\edb_top_inst/n2030 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/n2045 ), 
            .O(\edb_top_inst/n2046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3940 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3941  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8]), 
            .I1(\edb_top_inst/n1903 ), .I2(\edb_top_inst/n1906 ), .I3(\edb_top_inst/n2046 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3941 .LUTMASK = 16'hff80;
    EFX_LUT4 \edb_top_inst/LUT__3942  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), .I2(\edb_top_inst/la0/la_window_depth [1]), 
            .O(\edb_top_inst/n2047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3942 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3943  (.I0(\edb_top_inst/n2047 ), .I1(\edb_top_inst/n2043 ), 
            .I2(\edb_top_inst/la0/la_window_depth [0]), .O(\edb_top_inst/n2048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3943 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3944  (.I0(\edb_top_inst/n2048 ), .I1(\edb_top_inst/n2032 ), 
            .I2(\edb_top_inst/la0/la_window_depth [2]), .I3(\edb_top_inst/la0/la_window_depth [3]), 
            .O(\edb_top_inst/n2049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3944 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__3945  (.I0(\edb_top_inst/n2034 ), .I1(\edb_top_inst/la0/la_window_depth [2]), 
            .I2(\edb_top_inst/la0/la_window_depth [4]), .I3(\edb_top_inst/n2049 ), 
            .O(\edb_top_inst/n2050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3945 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3946  (.I0(\edb_top_inst/n1939 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9]), 
            .I2(\edb_top_inst/n2050 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3946 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3947  (.I0(\edb_top_inst/n1947 ), .I1(\edb_top_inst/n1906 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
            .I3(\edb_top_inst/n2018 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3947 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3948  (.I0(\edb_top_inst/n1895 ), .I1(\edb_top_inst/n1906 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1]), 
            .I3(\edb_top_inst/n2020 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3948 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3949  (.I0(\edb_top_inst/n1969 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2]), 
            .I2(\edb_top_inst/n2023 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3949 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3950  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3]), 
            .I1(\edb_top_inst/n2024 ), .I2(\edb_top_inst/n2027 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3950 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3951  (.I0(\edb_top_inst/n1900 ), .I1(\edb_top_inst/n2024 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4]), 
            .I3(\edb_top_inst/n2031 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3951 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3952  (.I0(\edb_top_inst/n1899 ), .I1(\edb_top_inst/n2024 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5]), 
            .I3(\edb_top_inst/n2035 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3952 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3953  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6]), 
            .I1(\edb_top_inst/n2036 ), .I2(\edb_top_inst/n2039 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3953 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3954  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/n1938 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7]), 
            .I3(\edb_top_inst/n2042 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3954 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3955  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8]), 
            .I1(\edb_top_inst/n1903 ), .I2(\edb_top_inst/n1906 ), .I3(\edb_top_inst/n2046 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3955 .LUTMASK = 16'hff80;
    EFX_LUT4 \edb_top_inst/LUT__3956  (.I0(\edb_top_inst/n1939 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9]), 
            .I2(\edb_top_inst/n2050 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3956 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3957  (.I0(\edb_top_inst/la0/opcode [0]), 
            .I1(\edb_top_inst/la0/opcode [3]), .I2(\edb_top_inst/la0/opcode [2]), 
            .I3(\edb_top_inst/la0/opcode [1]), .O(\edb_top_inst/la0/n594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3957 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3958  (.I0(\edb_top_inst/la0/module_state [1]), 
            .I1(\edb_top_inst/la0/module_state [2]), .I2(\edb_top_inst/la0/module_state [0]), 
            .I3(\edb_top_inst/la0/module_state [3]), .O(\edb_top_inst/n2051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3958 .LUTMASK = 16'hcc53;
    EFX_LUT4 \edb_top_inst/LUT__3959  (.I0(\edb_top_inst/n2051 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr [81]), .I3(jtag_inst1_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3959 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3960  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3960 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2993  (.I0(\edb_top_inst/la0/crc_data_out [24]), 
            .I1(\edb_top_inst/edb_user_dr [74]), .I2(\edb_top_inst/la0/crc_data_out [31]), 
            .I3(\edb_top_inst/edb_user_dr [81]), .O(\edb_top_inst/n1406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2993 .LUTMASK = 16'h9009;
    EFX_ADD \edb_top_inst/la0/add_417/i1  (.I0(\edb_top_inst/la0/address_counter [16]), 
            .I1(\edb_top_inst/la0/address_counter [15]), .CI(1'b0), .O(\edb_top_inst/la0/n1795 [1]), 
            .CO(\edb_top_inst/la0/add_417/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i1  (.I0(\edb_top_inst/la0/address_counter [0]), 
            .I1(\edb_top_inst/la0/n593 ), .CI(1'b0), .O(\edb_top_inst/la0/n1814 [0]), 
            .CO(\edb_top_inst/la0/add_98/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_419/i1  (.I0(\edb_top_inst/la0/bit_count [1]), 
            .I1(\edb_top_inst/la0/bit_count [0]), .CI(1'b0), .O(\edb_top_inst/la0/n1961 [1]), 
            .CO(\edb_top_inst/la0/add_419/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/add_419/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_419/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i1  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [1]), 
            .I1(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/trigger_skipper_n/n73 [1]), 
            .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(1'b1), .CI(n2336), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n342 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4660)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(1'b1), .CI(n2337), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n110 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4646)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10  (.I0(\edb_top_inst/la0/la_sample_cnt [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9  (.I0(\edb_top_inst/la0/la_sample_cnt [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [9]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8  (.I0(\edb_top_inst/la0/la_sample_cnt [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7  (.I0(\edb_top_inst/la0/la_sample_cnt [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6  (.I0(\edb_top_inst/la0/la_sample_cnt [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5  (.I0(\edb_top_inst/la0/la_sample_cnt [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4  (.I0(\edb_top_inst/la0/la_sample_cnt [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3  (.I0(\edb_top_inst/la0/la_sample_cnt [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n357 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [9]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n125 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer [0]), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n59 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4641)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), .CI(1'b0), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1  (.I0(\edb_top_inst/la0/la_sample_cnt [1]), 
            .I1(\edb_top_inst/la0/la_sample_cnt [0]), .CI(1'b0), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [1]), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt [0]), .CI(1'b0), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n22 [1]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4630)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [8]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [7]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [6]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [5]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [4]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [3]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n34 [2]), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4637)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i63  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [63]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n124 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i63 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i63 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i62  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [62]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n122 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [62]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i62 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i62 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i61  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [61]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n120 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [61]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i61 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i61 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i60  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [60]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n118 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [60]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i60 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i60 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i59  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [59]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n116 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [59]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i59 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i59 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i58  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [58]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n114 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [58]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i58 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i58 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i57  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [57]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n112 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [57]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i57 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i57 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i56  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [56]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n110 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [56]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i56 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i56 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i55  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [55]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n108 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [55]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i55 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i55 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i54  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [54]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n106 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [54]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i54 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i54 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i53  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [53]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n104 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [53]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i53 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i53 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i52  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [52]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n102 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [52]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i52 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i52 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i51  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [51]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n100 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [51]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i51 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i51 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i50  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [50]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n98 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [50]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i50 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i50 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i49  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [49]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n96 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [49]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i49 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i49 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i48  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [48]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n94 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [48]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i48 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i48 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i47  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [47]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n92 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [47]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i47 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i47 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i46  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [46]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n90 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [46]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i46 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i46 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i45  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [45]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n88 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [45]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i45 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i45 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i44  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [44]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n86 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [44]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i44 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i44 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i43  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [43]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n84 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [43]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i43 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i43 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i42  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [42]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n82 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [42]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i42 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i42 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i41  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [41]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n80 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [41]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i41 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i41 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i40  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [40]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n78 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [40]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i40 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i40 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i39  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [39]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n76 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [39]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i39 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i39 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i38  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [38]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n74 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [38]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i38 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i38 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i37  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [37]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n72 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [37]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i37 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i37 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i36  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [36]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n70 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [36]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i36 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i36 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i35  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [35]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n68 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [35]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i35 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i35 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i34  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [34]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n66 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [34]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i34 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i34 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i33  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [33]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n64 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [33]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i33 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i33 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i32  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [32]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n62 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [32]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i32 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i31  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [31]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n60 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [31]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i31 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i30  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [30]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n58 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [30]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i30 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i29  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [29]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n56 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [29]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i29 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i28  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [28]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n54 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [28]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i28 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i27  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [27]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n52 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [27]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i26  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [26]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n50 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [26]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i25  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [25]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n48 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [25]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i24  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n46 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [24]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i23  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n44 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [23]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i22  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n42 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [22]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i21  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n40 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [21]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i20  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n38 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [20]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i19  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n36 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [19]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i18  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n34 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [18]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i17  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n32 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [17]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i16  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [16]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n30 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [16]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i15  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [15]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n28 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [15]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i14  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [14]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n26 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [14]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i13  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [13]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n24 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [13]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i12  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [12]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n22 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [12]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i11  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [11]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n20 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [11]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i10  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n18 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [10]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i9  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n16 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [9]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i8  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n14 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [8]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i7  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n12 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [7]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i6  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n10 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [6]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i5  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n8 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [5]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i4  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n6 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [4]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i3  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n4 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [3]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/trigger_skipper_n/add_19/i2  (.I0(\edb_top_inst/la0/trigger_skipper_n/total_number_of_trigger_count [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/trigger_skipper_n/add_19/n2 ), 
            .O(\edb_top_inst/la0/trigger_skipper_n/n73 [2]), .CO(\edb_top_inst/la0/trigger_skipper_n/add_19/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(5830)
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/trigger_skipper_n/add_19/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_419/i5  (.I0(\edb_top_inst/la0/bit_count [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_419/n8 ), .O(\edb_top_inst/la0/n1961 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/add_419/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_419/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_419/i4  (.I0(\edb_top_inst/la0/bit_count [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_419/n6 ), .O(\edb_top_inst/la0/n1961 [4]), 
            .CO(\edb_top_inst/la0/add_419/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/add_419/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_419/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_419/i3  (.I0(\edb_top_inst/la0/bit_count [3]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_419/n4 ), .O(\edb_top_inst/la0/n1961 [3]), 
            .CO(\edb_top_inst/la0/add_419/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/add_419/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_419/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_419/i2  (.I0(\edb_top_inst/la0/bit_count [2]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_419/n2 ), .O(\edb_top_inst/la0/n1961 [2]), 
            .CO(\edb_top_inst/la0/add_419/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3697)
    defparam \edb_top_inst/la0/add_419/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_419/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i25  (.I0(\edb_top_inst/la0/address_counter [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n48 ), .O(\edb_top_inst/la0/n1814 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i24  (.I0(\edb_top_inst/la0/address_counter [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n46 ), .O(\edb_top_inst/la0/n1814 [23]), 
            .CO(\edb_top_inst/la0/add_98/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i23  (.I0(\edb_top_inst/la0/address_counter [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n44 ), .O(\edb_top_inst/la0/n1814 [22]), 
            .CO(\edb_top_inst/la0/add_98/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i22  (.I0(\edb_top_inst/la0/address_counter [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n42 ), .O(\edb_top_inst/la0/n1814 [21]), 
            .CO(\edb_top_inst/la0/add_98/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i21  (.I0(\edb_top_inst/la0/address_counter [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n40 ), .O(\edb_top_inst/la0/n1814 [20]), 
            .CO(\edb_top_inst/la0/add_98/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i20  (.I0(\edb_top_inst/la0/address_counter [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n38 ), .O(\edb_top_inst/la0/n1814 [19]), 
            .CO(\edb_top_inst/la0/add_98/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i19  (.I0(\edb_top_inst/la0/address_counter [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n36 ), .O(\edb_top_inst/la0/n1814 [18]), 
            .CO(\edb_top_inst/la0/add_98/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i18  (.I0(\edb_top_inst/la0/address_counter [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n34 ), .O(\edb_top_inst/la0/n1814 [17]), 
            .CO(\edb_top_inst/la0/add_98/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i17  (.I0(\edb_top_inst/la0/address_counter [16]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n32 ), .O(\edb_top_inst/la0/n1814 [16]), 
            .CO(\edb_top_inst/la0/add_98/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i16  (.I0(\edb_top_inst/la0/address_counter [15]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n30 ), .O(\edb_top_inst/la0/n1814 [15]), 
            .CO(\edb_top_inst/la0/add_98/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i15  (.I0(\edb_top_inst/la0/address_counter [14]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n28 ), .O(\edb_top_inst/la0/n1814 [14]), 
            .CO(\edb_top_inst/la0/add_98/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i14  (.I0(\edb_top_inst/la0/address_counter [13]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n26 ), .O(\edb_top_inst/la0/n1814 [13]), 
            .CO(\edb_top_inst/la0/add_98/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i13  (.I0(\edb_top_inst/la0/address_counter [12]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n24 ), .O(\edb_top_inst/la0/n1814 [12]), 
            .CO(\edb_top_inst/la0/add_98/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i12  (.I0(\edb_top_inst/la0/address_counter [11]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n22 ), .O(\edb_top_inst/la0/n1814 [11]), 
            .CO(\edb_top_inst/la0/add_98/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i11  (.I0(\edb_top_inst/la0/address_counter [10]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n20 ), .O(\edb_top_inst/la0/n1814 [10]), 
            .CO(\edb_top_inst/la0/add_98/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i10  (.I0(\edb_top_inst/la0/address_counter [9]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n18 ), .O(\edb_top_inst/la0/n1814 [9]), 
            .CO(\edb_top_inst/la0/add_98/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i9  (.I0(\edb_top_inst/la0/address_counter [8]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n16 ), .O(\edb_top_inst/la0/n1814 [8]), 
            .CO(\edb_top_inst/la0/add_98/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i8  (.I0(\edb_top_inst/la0/address_counter [7]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n14 ), .O(\edb_top_inst/la0/n1814 [7]), 
            .CO(\edb_top_inst/la0/add_98/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i7  (.I0(\edb_top_inst/la0/address_counter [6]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n12 ), .O(\edb_top_inst/la0/n1814 [6]), 
            .CO(\edb_top_inst/la0/add_98/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i6  (.I0(\edb_top_inst/la0/address_counter [5]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n10 ), .O(\edb_top_inst/la0/n1814 [5]), 
            .CO(\edb_top_inst/la0/add_98/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i5  (.I0(\edb_top_inst/la0/address_counter [4]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_98/n8 ), .O(\edb_top_inst/la0/n1814 [4]), 
            .CO(\edb_top_inst/la0/add_98/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i4  (.I0(\edb_top_inst/la0/address_counter [3]), 
            .I1(\edb_top_inst/la0/n596 ), .CI(\edb_top_inst/la0/add_98/n6 ), 
            .O(\edb_top_inst/la0/n1814 [3]), .CO(\edb_top_inst/la0/add_98/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i3  (.I0(\edb_top_inst/la0/address_counter [2]), 
            .I1(\edb_top_inst/la0/n595 ), .CI(\edb_top_inst/la0/add_98/n4 ), 
            .O(\edb_top_inst/la0/n1814 [2]), .CO(\edb_top_inst/la0/add_98/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_98/i2  (.I0(\edb_top_inst/la0/address_counter [1]), 
            .I1(\edb_top_inst/la0/n594 ), .CI(\edb_top_inst/la0/add_98/n2 ), 
            .O(\edb_top_inst/la0/n1814 [1]), .CO(\edb_top_inst/la0/add_98/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/add_98/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_98/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i9  (.I0(\edb_top_inst/la0/address_counter [24]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n16 ), .O(\edb_top_inst/la0/n1795 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i8  (.I0(\edb_top_inst/la0/address_counter [23]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n14 ), .O(\edb_top_inst/la0/n1795 [8]), 
            .CO(\edb_top_inst/la0/add_417/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i7  (.I0(\edb_top_inst/la0/address_counter [22]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n12 ), .O(\edb_top_inst/la0/n1795 [7]), 
            .CO(\edb_top_inst/la0/add_417/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i6  (.I0(\edb_top_inst/la0/address_counter [21]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n10 ), .O(\edb_top_inst/la0/n1795 [6]), 
            .CO(\edb_top_inst/la0/add_417/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i5  (.I0(\edb_top_inst/la0/address_counter [20]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n8 ), .O(\edb_top_inst/la0/n1795 [5]), 
            .CO(\edb_top_inst/la0/add_417/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i4  (.I0(\edb_top_inst/la0/address_counter [19]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n6 ), .O(\edb_top_inst/la0/n1795 [4]), 
            .CO(\edb_top_inst/la0/add_417/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i3  (.I0(\edb_top_inst/la0/address_counter [18]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n4 ), .O(\edb_top_inst/la0/n1795 [3]), 
            .CO(\edb_top_inst/la0/add_417/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_417/i2  (.I0(\edb_top_inst/la0/address_counter [17]), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_417/n2 ), .O(\edb_top_inst/la0/n1795 [2]), 
            .CO(\edb_top_inst/la0/add_417/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(3669)
    defparam \edb_top_inst/la0/add_417/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_417/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n576 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [9:5]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [9:5]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(406)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n576 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2 [4:0]}), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout [4:0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(406)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__6231 (.I0(b[0]), .I1(a[0]), .O(n30_2[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(36)
    defparam LUT__6231.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6232 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [4]), 
            .O(rx_data[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6232.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6233 (.I0(\uart_rx_inst/r_Clock_Count [3]), .I1(\uart_rx_inst/r_config_data [1]), 
            .I2(\uart_rx_inst/r_Clock_Count [0]), .I3(\uart_rx_inst/r_Clock_Count [1]), 
            .O(n2195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4ccf */ ;
    defparam LUT__6233.LUTMASK = 16'h4ccf;
    EFX_LUT4 LUT__6234 (.I0(\uart_rx_inst/r_config_data [1]), .I1(\uart_rx_inst/r_Clock_Count [6]), 
            .I2(\uart_rx_inst/r_Clock_Count [4]), .I3(\uart_rx_inst/r_Clock_Count [5]), 
            .O(n2196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__6234.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__6235 (.I0(n2195), .I1(n2196), .I2(\uart_rx_inst/r_Clock_Count [2]), 
            .O(n2197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6235.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6236 (.I0(\uart_rx_inst/r_Clock_Count [4]), .I1(\uart_rx_inst/r_Clock_Count [5]), 
            .O(n2198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6236.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6237 (.I0(\uart_rx_inst/r_Clock_Count [3]), .I1(n2198), 
            .I2(\uart_rx_inst/r_Clock_Count [6]), .I3(\uart_rx_inst/r_config_data [1]), 
            .O(n2199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__6237.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__6238 (.I0(n2199), .I1(n2197), .I2(\uart_rx_inst/r_Clock_Count [7]), 
            .I3(\uart_rx_inst/r_Clock_Count [8]), .O(n2200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6238.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6239 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(\uart_rx_inst/r_Clock_Count [29]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6239.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6240 (.I0(n2201), .I1(\uart_rx_inst/r_Clock_Count [26]), 
            .I2(\uart_rx_inst/r_Clock_Count [30]), .I3(\uart_rx_inst/r_config_data [1]), 
            .O(n2202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__6240.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__6241 (.I0(\uart_rx_inst/r_Clock_Count [24]), .I1(\uart_rx_inst/r_Clock_Count [25]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6241.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6242 (.I0(n2203), .I1(\uart_rx_inst/r_Clock_Count [20]), 
            .I2(\uart_rx_inst/r_Clock_Count [27]), .I3(\uart_rx_inst/r_config_data [1]), 
            .O(n2204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__6242.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__6243 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(\uart_rx_inst/r_Clock_Count [18]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6243.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6244 (.I0(\uart_rx_inst/r_Clock_Count [16]), .I1(\uart_rx_inst/r_Clock_Count [17]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6244.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6245 (.I0(\uart_rx_inst/r_Clock_Count [9]), .I1(\uart_rx_inst/r_Clock_Count [19]), 
            .I2(\uart_rx_inst/r_Clock_Count [31]), .I3(\uart_rx_inst/r_config_data [1]), 
            .O(n2207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6245.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6246 (.I0(\uart_rx_inst/r_Clock_Count [15]), .I1(\uart_rx_inst/r_Clock_Count [21]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6246.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6247 (.I0(n2205), .I1(n2206), .I2(n2207), .I3(n2208), 
            .O(n2209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6247.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6248 (.I0(\uart_rx_inst/r_Clock_Count [22]), .I1(\uart_rx_inst/r_Clock_Count [23]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6248.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6249 (.I0(\uart_rx_inst/r_Clock_Count [12]), .I1(\uart_rx_inst/r_Clock_Count [13]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6249.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6250 (.I0(\uart_rx_inst/r_Clock_Count [10]), .I1(\uart_rx_inst/r_Clock_Count [11]), 
            .I2(\uart_rx_inst/r_config_data [1]), .O(n2212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__6250.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__6251 (.I0(n2210), .I1(n2211), .I2(n2212), .O(n2213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6251.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6252 (.I0(n2202), .I1(n2204), .I2(n2209), .I3(n2213), 
            .O(n2214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6252.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6253 (.I0(\uart_rx_inst/r_SM_Main [2]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .O(\uart_rx_inst/n337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6253.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6254 (.I0(\uart_rx_inst/r_config_data [1]), .I1(n2200), 
            .I2(n2214), .I3(\uart_rx_inst/n337 ), .O(n2215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__6254.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__6255 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_Bit_Index [0]), 
            .O(n2216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6255.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6256 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(n2215), .I3(n2216), .O(\uart_rx_inst/n1220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6256.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6257 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [1]), .I3(\uart_rx_inst/r_Bit_Index [2]), 
            .O(n2217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6257.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6258 (.I0(\uart_rx_inst/r_SM_Main [1]), .I1(\uart_rx_inst/r_Rx_Data ), 
            .I2(\uart_rx_inst/r_SM_Main [0]), .O(n2218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6258.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6259 (.I0(\uart_rx_inst/r_config_data [1]), .I1(n2200), 
            .I2(n2214), .I3(\uart_rx_inst/r_SM_Main [1]), .O(n2219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__6259.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__6260 (.I0(n2205), .I1(n2206), .O(n2220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6260.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6261 (.I0(n2210), .I1(n2211), .O(n2221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6261.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6262 (.I0(\uart_rx_inst/r_Clock_Count [6]), .I1(\uart_rx_inst/r_Clock_Count [7]), 
            .O(n2222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6262.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6263 (.I0(\uart_rx_inst/r_Clock_Count [31]), .I1(\uart_rx_inst/r_Clock_Count [3]), 
            .I2(\uart_rx_inst/r_Clock_Count [4]), .I3(\uart_rx_inst/r_Clock_Count [1]), 
            .O(n2223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6263.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6264 (.I0(n2222), .I1(n2223), .O(n2224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6264.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6265 (.I0(n2202), .I1(n2220), .I2(n2221), .I3(n2224), 
            .O(n2225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6265.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6266 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [2]), 
            .I2(\uart_rx_inst/r_Clock_Count [5]), .I3(\uart_rx_inst/r_Clock_Count [8]), 
            .O(n2226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6266.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6267 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [9]), 
            .I2(\uart_rx_inst/r_Clock_Count [19]), .I3(\uart_rx_inst/r_config_data [1]), 
            .O(n2227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6267.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6268 (.I0(n2212), .I1(\uart_rx_inst/r_Clock_Count [21]), 
            .I2(\uart_rx_inst/r_Clock_Count [15]), .I3(\uart_rx_inst/r_Clock_Count [10]), 
            .O(n2228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__6268.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__6269 (.I0(n2226), .I1(n2227), .I2(n2204), .I3(n2228), 
            .O(n2229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6269.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6270 (.I0(n2229), .I1(n2225), .I2(\uart_rx_inst/r_SM_Main [1]), 
            .I3(\uart_rx_inst/r_SM_Main [0]), .O(n2230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6270.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6271 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n2230), 
            .O(\uart_rx_inst/n1145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf03b */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6271.LUTMASK = 16'hf03b;
    EFX_LUT4 LUT__6272 (.I0(n2229), .I1(n2225), .I2(\uart_rx_inst/r_SM_Main [1]), 
            .I3(\uart_rx_inst/r_SM_Main [0]), .O(n2231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6272.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6273 (.I0(n2231), .I1(n2219), .I2(\uart_rx_inst/r_Clock_Count [0]), 
            .O(\uart_rx_inst/n1148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6273.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6274 (.I0(n2225), .I1(n2229), .O(n2232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6274.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6275 (.I0(\uart_rx_inst/r_Rx_Data ), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(\uart_rx_inst/r_SM_Main [0]), .O(n2233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6275.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6276 (.I0(n2233), .I1(n2232), .I2(\uart_rx_inst/r_SM_Main [2]), 
            .O(ceg_net14)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(80)
    defparam LUT__6276.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__6277 (.I0(\uart_rx_inst/r_config_data [1]), .I1(n2200), 
            .I2(n2214), .O(\uart_rx_inst/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(129)
    defparam LUT__6277.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6278 (.I0(\uart_rx_inst/n151 ), .I1(\uart_rx_inst/r_SM_Main [2]), 
            .I2(\uart_rx_inst/r_SM_Main [1]), .I3(\uart_rx_inst/r_SM_Main [0]), 
            .O(ceg_net32)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(80)
    defparam LUT__6278.LUTMASK = 16'heff0;
    EFX_LUT4 LUT__6279 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .O(\uart_rx_inst/n1152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(143)
    defparam LUT__6279.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6280 (.I0(n2219), .I1(\uart_rx_inst/r_SM_Main [0]), .I2(\uart_rx_inst/r_SM_Main [2]), 
            .O(ceg_net26)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(80)
    defparam LUT__6280.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__6281 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_Bit_Index [0]), 
            .O(n2234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6281.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6282 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(n2215), .I3(n2234), .O(\uart_rx_inst/n1199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6282.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6283 (.I0(\uart_rx_inst/n337 ), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .O(n2235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6283.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6284 (.I0(\uart_rx_inst/n151 ), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(n2216), .I3(n2235), .O(\uart_rx_inst/n1202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6284.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6285 (.I0(\uart_rx_inst/n151 ), .I1(\uart_rx_inst/r_Bit_Index [2]), 
            .I2(n2234), .I3(n2235), .O(\uart_rx_inst/n1205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6285.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6286 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(n2216), 
            .I2(n2215), .I3(\uart_rx_inst/r_Bit_Index [2]), .O(\uart_rx_inst/n1208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6286.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6287 (.I0(\uart_rx_inst/r_Bit_Index [1]), .I1(n2234), 
            .I2(n2215), .I3(\uart_rx_inst/r_Bit_Index [2]), .O(\uart_rx_inst/n1211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6287.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6288 (.I0(\uart_rx_inst/n151 ), .I1(n2235), .I2(n2216), 
            .I3(\uart_rx_inst/r_Bit_Index [2]), .O(\uart_rx_inst/n1214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6288.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6289 (.I0(\uart_rx_inst/n151 ), .I1(n2235), .I2(n2234), 
            .I3(\uart_rx_inst/r_Bit_Index [2]), .O(\uart_rx_inst/n1217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6289.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6290 (.I0(\uart_rx_inst/r_Rx_Data ), .I1(\uart_rx_inst/r_SM_Main [0]), 
            .O(n2236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6290.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6291 (.I0(\uart_rx_inst/r_config_data [1]), .I1(n2200), 
            .I2(n2214), .I3(\uart_rx_inst/r_SM_Main [0]), .O(n2237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__6291.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__6292 (.I0(n2236), .I1(n2232), .I2(\uart_rx_inst/r_SM_Main [1]), 
            .I3(n2237), .O(\uart_rx_inst/n826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6292.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__6293 (.I0(\uart_rx_inst/n337 ), .I1(\uart_rx_inst/r_SM_Main [0]), 
            .O(\uart_rx_inst/n1180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6293.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6294 (.I0(n2219), .I1(n2231), .I2(\uart_rx_inst/r_Clock_Count [0]), 
            .I3(\uart_rx_inst/r_Clock_Count [1]), .O(\uart_rx_inst/n833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6294.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6295 (.I0(\uart_rx_inst/r_Clock_Count [0]), .I1(\uart_rx_inst/r_Clock_Count [1]), 
            .O(n2238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6295.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6296 (.I0(n2219), .I1(n2231), .I2(n2238), .I3(\uart_rx_inst/r_Clock_Count [2]), 
            .O(\uart_rx_inst/n836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6296.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6297 (.I0(n2238), .I1(\uart_rx_inst/r_Clock_Count [2]), 
            .I2(\uart_rx_inst/r_Clock_Count [3]), .O(n2239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6297.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6298 (.I0(n2231), .I1(n2219), .I2(n2239), .O(\uart_rx_inst/n839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6298.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6299 (.I0(n2238), .I1(\uart_rx_inst/r_Clock_Count [2]), 
            .I2(\uart_rx_inst/r_Clock_Count [3]), .O(n2240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6299.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6300 (.I0(n2219), .I1(n2231), .I2(n2240), .I3(\uart_rx_inst/r_Clock_Count [4]), 
            .O(\uart_rx_inst/n842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6300.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6301 (.I0(n2240), .I1(\uart_rx_inst/r_Clock_Count [4]), 
            .I2(\uart_rx_inst/r_Clock_Count [5]), .O(n2241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6301.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6302 (.I0(n2231), .I1(n2219), .I2(n2241), .O(\uart_rx_inst/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6302.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6303 (.I0(n2198), .I1(n2238), .I2(\uart_rx_inst/r_Clock_Count [2]), 
            .I3(\uart_rx_inst/r_Clock_Count [3]), .O(n2242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6303.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6304 (.I0(n2219), .I1(n2231), .I2(n2242), .I3(\uart_rx_inst/r_Clock_Count [6]), 
            .O(\uart_rx_inst/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6304.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6305 (.I0(n2242), .I1(\uart_rx_inst/r_Clock_Count [6]), 
            .I2(\uart_rx_inst/r_Clock_Count [7]), .O(n2243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6305.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6306 (.I0(n2231), .I1(n2219), .I2(n2243), .O(\uart_rx_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6306.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6307 (.I0(n2242), .I1(n2222), .O(n2244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6307.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6308 (.I0(n2219), .I1(n2231), .I2(n2244), .I3(\uart_rx_inst/r_Clock_Count [8]), 
            .O(\uart_rx_inst/n854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6308.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6309 (.I0(n2244), .I1(\uart_rx_inst/r_Clock_Count [8]), 
            .I2(\uart_rx_inst/r_Clock_Count [9]), .O(n2245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6309.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6310 (.I0(n2231), .I1(n2219), .I2(n2245), .O(\uart_rx_inst/n857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6310.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6311 (.I0(\uart_rx_inst/r_Clock_Count [8]), .I1(\uart_rx_inst/r_Clock_Count [9]), 
            .O(n2246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6311.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6312 (.I0(n2244), .I1(n2246), .I2(\uart_rx_inst/r_Clock_Count [10]), 
            .O(n2247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6312.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6313 (.I0(n2231), .I1(n2219), .I2(n2247), .O(\uart_rx_inst/n860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6313.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6314 (.I0(n2242), .I1(n2246), .O(n2248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6314.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6315 (.I0(n2248), .I1(n2222), .I2(\uart_rx_inst/r_Clock_Count [10]), 
            .O(n2249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6315.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6316 (.I0(n2219), .I1(n2231), .I2(n2249), .I3(\uart_rx_inst/r_Clock_Count [11]), 
            .O(\uart_rx_inst/n863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6316.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6317 (.I0(\uart_rx_inst/r_Clock_Count [6]), .I1(\uart_rx_inst/r_Clock_Count [7]), 
            .I2(\uart_rx_inst/r_Clock_Count [10]), .I3(\uart_rx_inst/r_Clock_Count [11]), 
            .O(n2250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6317.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6318 (.I0(n2248), .I1(n2250), .O(n2251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6318.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6319 (.I0(n2219), .I1(n2231), .I2(n2251), .I3(\uart_rx_inst/r_Clock_Count [12]), 
            .O(\uart_rx_inst/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6319.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6320 (.I0(n2248), .I1(n2250), .I2(\uart_rx_inst/r_Clock_Count [12]), 
            .I3(\uart_rx_inst/r_Clock_Count [13]), .O(n2252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6320.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6321 (.I0(n2231), .I1(n2219), .I2(n2252), .O(\uart_rx_inst/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6321.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6322 (.I0(n2246), .I1(n2250), .I2(\uart_rx_inst/r_Clock_Count [12]), 
            .I3(\uart_rx_inst/r_Clock_Count [13]), .O(n2253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6322.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6323 (.I0(n2242), .I1(n2253), .I2(\uart_rx_inst/r_Clock_Count [14]), 
            .O(n2254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6323.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6324 (.I0(n2231), .I1(n2219), .I2(n2254), .O(\uart_rx_inst/n872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6324.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6325 (.I0(n2242), .I1(n2253), .I2(\uart_rx_inst/r_Clock_Count [14]), 
            .I3(\uart_rx_inst/r_Clock_Count [15]), .O(n2255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6325.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6326 (.I0(n2231), .I1(n2219), .I2(n2255), .O(\uart_rx_inst/n875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6326.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6327 (.I0(n2242), .I1(\uart_rx_inst/r_Clock_Count [14]), 
            .I2(\uart_rx_inst/r_Clock_Count [15]), .O(n2256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6327.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6328 (.I0(n2256), .I1(n2253), .O(n2257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6328.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6329 (.I0(n2219), .I1(n2231), .I2(n2257), .I3(\uart_rx_inst/r_Clock_Count [16]), 
            .O(\uart_rx_inst/n878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6329.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6330 (.I0(n2256), .I1(n2253), .I2(\uart_rx_inst/r_Clock_Count [16]), 
            .I3(\uart_rx_inst/r_Clock_Count [17]), .O(n2258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6330.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6331 (.I0(n2231), .I1(n2219), .I2(n2258), .O(\uart_rx_inst/n881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6331.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6332 (.I0(n2242), .I1(n2246), .I2(\uart_rx_inst/r_Clock_Count [14]), 
            .I3(\uart_rx_inst/r_Clock_Count [15]), .O(n2259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6332.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6333 (.I0(n2250), .I1(\uart_rx_inst/r_Clock_Count [12]), 
            .I2(\uart_rx_inst/r_Clock_Count [13]), .O(n2260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6333.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6334 (.I0(n2260), .I1(\uart_rx_inst/r_Clock_Count [16]), 
            .I2(\uart_rx_inst/r_Clock_Count [17]), .O(n2261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6334.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6335 (.I0(n2259), .I1(n2261), .I2(\uart_rx_inst/r_Clock_Count [18]), 
            .O(n2262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6335.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6336 (.I0(n2231), .I1(n2219), .I2(n2262), .O(\uart_rx_inst/n884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6336.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6337 (.I0(n2259), .I1(n2261), .I2(\uart_rx_inst/r_Clock_Count [18]), 
            .I3(\uart_rx_inst/r_Clock_Count [19]), .O(n2263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6337.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6338 (.I0(n2231), .I1(n2219), .I2(n2263), .O(\uart_rx_inst/n887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6338.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6339 (.I0(\uart_rx_inst/r_Clock_Count [14]), .I1(\uart_rx_inst/r_Clock_Count [15]), 
            .I2(\uart_rx_inst/r_Clock_Count [18]), .I3(\uart_rx_inst/r_Clock_Count [19]), 
            .O(n2264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6339.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6340 (.I0(n2248), .I1(n2261), .I2(n2264), .O(n2265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6340.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6341 (.I0(n2219), .I1(n2231), .I2(n2265), .I3(\uart_rx_inst/r_Clock_Count [20]), 
            .O(\uart_rx_inst/n890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6341.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6342 (.I0(n2248), .I1(n2261), .I2(n2264), .I3(\uart_rx_inst/r_Clock_Count [20]), 
            .O(n2266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6342.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6343 (.I0(n2219), .I1(n2231), .I2(n2266), .I3(\uart_rx_inst/r_Clock_Count [21]), 
            .O(\uart_rx_inst/n893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6343.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6344 (.I0(n2242), .I1(n2264), .I2(\uart_rx_inst/r_Clock_Count [12]), 
            .I3(\uart_rx_inst/r_Clock_Count [13]), .O(n2267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6344.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6345 (.I0(\uart_rx_inst/r_Clock_Count [16]), .I1(\uart_rx_inst/r_Clock_Count [17]), 
            .I2(\uart_rx_inst/r_Clock_Count [20]), .I3(\uart_rx_inst/r_Clock_Count [21]), 
            .O(n2268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6345.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6346 (.I0(n2246), .I1(n2250), .I2(n2268), .O(n2269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6346.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6347 (.I0(n2267), .I1(n2269), .O(n2270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6347.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6348 (.I0(n2219), .I1(n2231), .I2(n2270), .I3(\uart_rx_inst/r_Clock_Count [22]), 
            .O(\uart_rx_inst/n896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6348.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6349 (.I0(n2267), .I1(n2269), .I2(\uart_rx_inst/r_Clock_Count [22]), 
            .O(n2271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6349.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6350 (.I0(n2219), .I1(n2231), .I2(n2271), .I3(\uart_rx_inst/r_Clock_Count [23]), 
            .O(\uart_rx_inst/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6350.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6351 (.I0(n2246), .I1(n2268), .I2(\uart_rx_inst/r_Clock_Count [22]), 
            .I3(\uart_rx_inst/r_Clock_Count [23]), .O(n2272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6351.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6352 (.I0(n2242), .I1(n2260), .I2(n2272), .I3(n2264), 
            .O(n2273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6352.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6353 (.I0(n2219), .I1(n2231), .I2(n2273), .I3(\uart_rx_inst/r_Clock_Count [24]), 
            .O(\uart_rx_inst/n902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6353.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6354 (.I0(n2273), .I1(\uart_rx_inst/r_Clock_Count [24]), 
            .I2(\uart_rx_inst/r_Clock_Count [25]), .O(n2274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6354.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6355 (.I0(n2231), .I1(n2219), .I2(n2274), .O(\uart_rx_inst/n905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6355.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6356 (.I0(n2198), .I1(n2264), .I2(\uart_rx_inst/r_Clock_Count [24]), 
            .I3(\uart_rx_inst/r_Clock_Count [25]), .O(n2275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6356.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6357 (.I0(n2240), .I1(n2253), .I2(n2275), .I3(n2272), 
            .O(n2276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6357.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6358 (.I0(n2219), .I1(n2231), .I2(n2276), .I3(\uart_rx_inst/r_Clock_Count [26]), 
            .O(\uart_rx_inst/n908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6358.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6359 (.I0(n2276), .I1(\uart_rx_inst/r_Clock_Count [26]), 
            .I2(\uart_rx_inst/r_Clock_Count [27]), .O(n2277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6359.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6360 (.I0(n2231), .I1(n2219), .I2(n2277), .O(\uart_rx_inst/n911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6360.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6361 (.I0(\uart_rx_inst/r_Clock_Count [24]), .I1(\uart_rx_inst/r_Clock_Count [25]), 
            .I2(\uart_rx_inst/r_Clock_Count [26]), .I3(\uart_rx_inst/r_Clock_Count [27]), 
            .O(n2278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6361.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6362 (.I0(n2272), .I1(n2222), .I2(n2278), .O(n2279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6362.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6363 (.I0(\uart_rx_inst/r_Clock_Count [10]), .I1(\uart_rx_inst/r_Clock_Count [11]), 
            .O(n2280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6363.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6364 (.I0(n2267), .I1(n2279), .I2(n2280), .O(n2281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6364.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6365 (.I0(n2219), .I1(n2231), .I2(n2281), .I3(\uart_rx_inst/r_Clock_Count [28]), 
            .O(\uart_rx_inst/n914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6365.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6366 (.I0(n2267), .I1(n2279), .I2(n2280), .I3(\uart_rx_inst/r_Clock_Count [28]), 
            .O(n2282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6366.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6367 (.I0(n2219), .I1(n2231), .I2(n2282), .I3(\uart_rx_inst/r_Clock_Count [29]), 
            .O(\uart_rx_inst/n917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6367.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6368 (.I0(\uart_rx_inst/r_Clock_Count [28]), .I1(\uart_rx_inst/r_Clock_Count [29]), 
            .O(n2283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6368.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6369 (.I0(n2267), .I1(n2279), .I2(n2283), .I3(n2280), 
            .O(n2284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6369.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6370 (.I0(n2219), .I1(n2231), .I2(n2284), .I3(\uart_rx_inst/r_Clock_Count [30]), 
            .O(\uart_rx_inst/n920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6370.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6371 (.I0(n2283), .I1(\uart_rx_inst/r_Clock_Count [30]), 
            .O(n2285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6371.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6372 (.I0(n2267), .I1(n2279), .I2(n2285), .I3(n2280), 
            .O(n2286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6372.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6373 (.I0(n2219), .I1(n2231), .I2(n2286), .I3(\uart_rx_inst/r_Clock_Count [31]), 
            .O(\uart_rx_inst/n923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ee0 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(167)
    defparam LUT__6373.LUTMASK = 16'h0ee0;
    EFX_LUT4 LUT__6374 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_SM_Main [1]), .O(\uart_rx_inst/n927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(143)
    defparam LUT__6374.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6375 (.I0(\uart_rx_inst/r_Bit_Index [0]), .I1(\uart_rx_inst/r_Bit_Index [1]), 
            .I2(\uart_rx_inst/r_Bit_Index [2]), .I3(\uart_rx_inst/r_SM_Main [1]), 
            .O(\uart_rx_inst/n931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(143)
    defparam LUT__6375.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6376 (.I0(\uart_rx_inst/r_SM_Main [0]), .I1(\uart_rx_inst/r_SM_Main [1]), 
            .I2(\uart_rx_inst/r_SM_Main [2]), .O(\uart_rx_inst/n1161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(17)
    defparam LUT__6376.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__6377 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [1]), 
            .O(rx_data[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6377.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6378 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [2]), 
            .O(rx_data[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6378.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6379 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [3]), 
            .O(rx_data[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6379.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6380 (.I0(b[1]), .I1(a[1]), .O(n25[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(35)
    defparam LUT__6380.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6381 (.I0(b[2]), .I1(a[2]), .O(n25[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(35)
    defparam LUT__6381.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6382 (.I0(b[3]), .I1(a[3]), .O(n25[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(35)
    defparam LUT__6382.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6383 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_config_data [31]), 
            .I2(\uart_tx_inst/r_Clock_Count [1]), .I3(\uart_tx_inst/r_Clock_Count [2]), 
            .O(n2287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__6383.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__6384 (.I0(\uart_tx_inst/r_Clock_Count [4]), .I1(\uart_tx_inst/r_Clock_Count [5]), 
            .O(n2288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6384.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6385 (.I0(n2287), .I1(\uart_tx_inst/r_config_data [31]), 
            .I2(\uart_tx_inst/r_Clock_Count [3]), .I3(n2288), .O(n2289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__6385.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__6386 (.I0(\uart_tx_inst/r_Clock_Count [7]), .I1(\uart_tx_inst/r_Clock_Count [8]), 
            .O(n2290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6386.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6387 (.I0(n2289), .I1(\uart_tx_inst/r_config_data [31]), 
            .I2(\uart_tx_inst/r_Clock_Count [6]), .I3(n2290), .O(n2291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__6387.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__6388 (.I0(\uart_tx_inst/r_SM_Main [0]), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .O(n2292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6388.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6389 (.I0(\uart_tx_inst/r_Clock_Count [10]), .I1(\uart_tx_inst/r_Clock_Count [11]), 
            .I2(\uart_tx_inst/r_Clock_Count [14]), .I3(\uart_tx_inst/r_Clock_Count [15]), 
            .O(n2293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6389.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6390 (.I0(n2293), .I1(\uart_tx_inst/r_Clock_Count [24]), 
            .I2(\uart_tx_inst/r_Clock_Count [25]), .I3(\uart_tx_inst/r_Clock_Count [10]), 
            .O(n2294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__6390.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__6391 (.I0(\uart_tx_inst/r_Clock_Count [10]), .I1(\uart_tx_inst/r_Clock_Count [27]), 
            .I2(\uart_tx_inst/r_Clock_Count [30]), .I3(\uart_tx_inst/r_config_data [31]), 
            .O(n2295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6391.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6392 (.I0(\uart_tx_inst/r_Clock_Count [9]), .I1(\uart_tx_inst/r_Clock_Count [12]), 
            .I2(\uart_tx_inst/r_Clock_Count [13]), .I3(\uart_tx_inst/r_Clock_Count [16]), 
            .O(n2296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6392.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6393 (.I0(\uart_tx_inst/r_Clock_Count [10]), .I1(\uart_tx_inst/r_Clock_Count [18]), 
            .I2(\uart_tx_inst/r_Clock_Count [19]), .I3(\uart_tx_inst/r_Clock_Count [26]), 
            .O(n2297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6393.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6394 (.I0(\uart_tx_inst/r_Clock_Count [9]), .I1(\uart_tx_inst/r_Clock_Count [17]), 
            .I2(\uart_tx_inst/r_Clock_Count [20]), .I3(\uart_tx_inst/r_Clock_Count [21]), 
            .O(n2298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6394.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6395 (.I0(\uart_tx_inst/r_Clock_Count [9]), .I1(\uart_tx_inst/r_Clock_Count [22]), 
            .I2(\uart_tx_inst/r_Clock_Count [23]), .I3(\uart_tx_inst/r_Clock_Count [28]), 
            .O(n2299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6395.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6396 (.I0(\uart_tx_inst/r_Clock_Count [9]), .I1(\uart_tx_inst/r_Clock_Count [29]), 
            .I2(\uart_tx_inst/r_Clock_Count [31]), .I3(\uart_tx_inst/r_config_data [31]), 
            .O(n2300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__6396.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__6397 (.I0(n2297), .I1(n2298), .I2(n2299), .I3(n2300), 
            .O(n2301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6397.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6398 (.I0(n2295), .I1(n2296), .I2(n2294), .I3(n2301), 
            .O(n2302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6398.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6399 (.I0(\uart_tx_inst/r_config_data [31]), .I1(n2291), 
            .I2(n2292), .I3(n2302), .O(n2303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__6399.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__6400 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(n2303), 
            .O(\uart_tx_inst/n1116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6400.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6401 (.I0(\uart_tx_inst/r_Tx_Data [4]), .I1(\uart_tx_inst/r_Tx_Data [6]), 
            .I2(\uart_tx_inst/r_Bit_Index [0]), .I3(\uart_tx_inst/r_Bit_Index [1]), 
            .O(n2304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6401.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6402 (.I0(\uart_tx_inst/r_Tx_Data [5]), .I1(\uart_tx_inst/r_Tx_Data [7]), 
            .I2(\uart_tx_inst/r_Bit_Index [1]), .I3(\uart_tx_inst/r_Bit_Index [0]), 
            .O(n2305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6402.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6403 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_Tx_Data [3]), .O(n2306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6403.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6404 (.I0(n2305), .I1(n2304), .I2(n2306), .I3(\uart_tx_inst/r_Bit_Index [2]), 
            .O(n2307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__6404.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__6405 (.I0(n2307), .I1(\uart_tx_inst/r_SM_Main [0]), .I2(\uart_tx_inst/r_SM_Main [1]), 
            .O(\uart_tx_inst/n733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(287)
    defparam LUT__6405.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6406 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .O(\uart_tx_inst/n1120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(260)
    defparam LUT__6406.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6407 (.I0(\uart_tx_inst/r_config_data [31]), .I1(n2291), 
            .I2(n2302), .O(\uart_tx_inst/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(234)
    defparam LUT__6407.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6408 (.I0(\uart_tx_inst/r_SM_Main [1]), .I1(\uart_tx_inst/n50 ), 
            .I2(\uart_tx_inst/r_SM_Main [0]), .I3(\uart_tx_inst/r_SM_Main [2]), 
            .O(ceg_net28)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(203)
    defparam LUT__6408.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__6409 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_Bit_Index [2]), .I3(\uart_tx_inst/r_SM_Main [1]), 
            .O(n2308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6409.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6410 (.I0(\uart_tx_inst/r_SM_Main [1]), .I1(send), .O(n2309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6410.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6411 (.I0(n2308), .I1(n2309), .I2(\uart_tx_inst/n50 ), 
            .I3(\uart_tx_inst/r_SM_Main [0]), .O(\uart_tx_inst/n1112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ce */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(287)
    defparam LUT__6411.LUTMASK = 16'hf0ce;
    EFX_LUT4 LUT__6412 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(n2303), .O(\uart_tx_inst/n786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6412.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6413 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(\uart_tx_inst/r_Clock_Count [2]), .I3(n2303), .O(\uart_tx_inst/n789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6413.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6414 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(\uart_tx_inst/r_Clock_Count [2]), .I3(\uart_tx_inst/r_Clock_Count [3]), 
            .O(n2310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6414.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6415 (.I0(n2310), .I1(n2303), .O(\uart_tx_inst/n792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6415.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6416 (.I0(\uart_tx_inst/r_Clock_Count [0]), .I1(\uart_tx_inst/r_Clock_Count [1]), 
            .I2(\uart_tx_inst/r_Clock_Count [2]), .I3(\uart_tx_inst/r_Clock_Count [3]), 
            .O(n2311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6416.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6417 (.I0(n2311), .I1(\uart_tx_inst/r_Clock_Count [4]), 
            .I2(n2303), .O(\uart_tx_inst/n795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6417.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6418 (.I0(n2311), .I1(\uart_tx_inst/r_Clock_Count [4]), 
            .I2(\uart_tx_inst/r_Clock_Count [5]), .I3(n2303), .O(\uart_tx_inst/n798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6418.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6419 (.I0(n2288), .I1(n2311), .O(n2312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6419.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6420 (.I0(n2312), .I1(\uart_tx_inst/r_Clock_Count [6]), 
            .I2(n2303), .O(\uart_tx_inst/n801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6420.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6421 (.I0(n2312), .I1(\uart_tx_inst/r_Clock_Count [6]), 
            .I2(\uart_tx_inst/r_Clock_Count [7]), .I3(n2303), .O(\uart_tx_inst/n804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6421.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6422 (.I0(n2312), .I1(\uart_tx_inst/r_Clock_Count [6]), 
            .I2(\uart_tx_inst/r_Clock_Count [7]), .O(n2313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6422.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6423 (.I0(n2313), .I1(\uart_tx_inst/r_Clock_Count [8]), 
            .I2(n2303), .O(\uart_tx_inst/n807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6423.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6424 (.I0(n2313), .I1(\uart_tx_inst/r_Clock_Count [8]), 
            .I2(\uart_tx_inst/r_Clock_Count [9]), .I3(n2303), .O(\uart_tx_inst/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6424.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6425 (.I0(n2313), .I1(\uart_tx_inst/r_Clock_Count [8]), 
            .I2(\uart_tx_inst/r_Clock_Count [9]), .O(n2314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6425.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6426 (.I0(n2314), .I1(\uart_tx_inst/r_Clock_Count [10]), 
            .I2(n2303), .O(\uart_tx_inst/n813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6426.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6427 (.I0(n2314), .I1(\uart_tx_inst/r_Clock_Count [10]), 
            .I2(\uart_tx_inst/r_Clock_Count [11]), .I3(n2303), .O(\uart_tx_inst/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6427.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6428 (.I0(\uart_tx_inst/r_Clock_Count [8]), .I1(\uart_tx_inst/r_Clock_Count [9]), 
            .I2(\uart_tx_inst/r_Clock_Count [10]), .I3(\uart_tx_inst/r_Clock_Count [11]), 
            .O(n2315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6428.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6429 (.I0(n2312), .I1(n2315), .I2(\uart_tx_inst/r_Clock_Count [6]), 
            .I3(\uart_tx_inst/r_Clock_Count [7]), .O(n2316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6429.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6430 (.I0(n2316), .I1(\uart_tx_inst/r_Clock_Count [12]), 
            .I2(n2303), .O(\uart_tx_inst/n819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6430.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6431 (.I0(n2316), .I1(\uart_tx_inst/r_Clock_Count [12]), 
            .I2(\uart_tx_inst/r_Clock_Count [13]), .I3(n2303), .O(\uart_tx_inst/n822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6431.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6432 (.I0(\uart_tx_inst/r_Clock_Count [6]), .I1(\uart_tx_inst/r_Clock_Count [7]), 
            .I2(\uart_tx_inst/r_Clock_Count [12]), .I3(\uart_tx_inst/r_Clock_Count [13]), 
            .O(n2317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6432.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6433 (.I0(n2312), .I1(n2315), .I2(n2317), .O(n2318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6433.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6434 (.I0(n2318), .I1(\uart_tx_inst/r_Clock_Count [14]), 
            .I2(n2303), .O(\uart_tx_inst/n825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6434.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6435 (.I0(n2318), .I1(\uart_tx_inst/r_Clock_Count [14]), 
            .I2(\uart_tx_inst/r_Clock_Count [15]), .I3(n2303), .O(\uart_tx_inst/n828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6435.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6436 (.I0(n2318), .I1(\uart_tx_inst/r_Clock_Count [14]), 
            .I2(\uart_tx_inst/r_Clock_Count [15]), .O(n2319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6436.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6437 (.I0(n2319), .I1(\uart_tx_inst/r_Clock_Count [16]), 
            .I2(n2303), .O(\uart_tx_inst/n831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6437.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6438 (.I0(n2319), .I1(\uart_tx_inst/r_Clock_Count [16]), 
            .I2(\uart_tx_inst/r_Clock_Count [17]), .I3(n2303), .O(\uart_tx_inst/n834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6438.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6439 (.I0(\uart_tx_inst/r_Clock_Count [14]), .I1(\uart_tx_inst/r_Clock_Count [15]), 
            .I2(\uart_tx_inst/r_Clock_Count [16]), .I3(\uart_tx_inst/r_Clock_Count [17]), 
            .O(n2320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6439.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6440 (.I0(n2318), .I1(n2320), .O(n2321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6440.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6441 (.I0(n2321), .I1(\uart_tx_inst/r_Clock_Count [18]), 
            .I2(n2303), .O(\uart_tx_inst/n837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6441.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6442 (.I0(n2321), .I1(\uart_tx_inst/r_Clock_Count [18]), 
            .I2(\uart_tx_inst/r_Clock_Count [19]), .I3(n2303), .O(\uart_tx_inst/n840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6442.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6443 (.I0(\uart_tx_inst/r_Clock_Count [18]), .I1(\uart_tx_inst/r_Clock_Count [19]), 
            .O(n2322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6443.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6444 (.I0(n2321), .I1(n2322), .I2(\uart_tx_inst/r_Clock_Count [20]), 
            .I3(n2303), .O(\uart_tx_inst/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6444.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6445 (.I0(n2318), .I1(n2322), .I2(n2320), .I3(\uart_tx_inst/r_Clock_Count [20]), 
            .O(n2323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6445.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6446 (.I0(n2323), .I1(\uart_tx_inst/r_Clock_Count [21]), 
            .I2(n2303), .O(\uart_tx_inst/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6446.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6447 (.I0(n2322), .I1(\uart_tx_inst/r_Clock_Count [20]), 
            .I2(\uart_tx_inst/r_Clock_Count [21]), .O(n2324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6447.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6448 (.I0(n2318), .I1(n2324), .I2(n2320), .O(n2325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6448.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6449 (.I0(n2325), .I1(\uart_tx_inst/r_Clock_Count [22]), 
            .I2(n2303), .O(\uart_tx_inst/n849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6449.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6450 (.I0(n2325), .I1(\uart_tx_inst/r_Clock_Count [22]), 
            .I2(\uart_tx_inst/r_Clock_Count [23]), .I3(n2303), .O(\uart_tx_inst/n852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6450.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6451 (.I0(\uart_tx_inst/r_Clock_Count [22]), .I1(\uart_tx_inst/r_Clock_Count [23]), 
            .O(n2326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6451.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6452 (.I0(n2325), .I1(n2326), .I2(\uart_tx_inst/r_Clock_Count [24]), 
            .I3(n2303), .O(\uart_tx_inst/n855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6452.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6453 (.I0(n2326), .I1(\uart_tx_inst/r_Clock_Count [24]), 
            .O(n2327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6453.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6454 (.I0(n2325), .I1(n2327), .I2(\uart_tx_inst/r_Clock_Count [25]), 
            .I3(n2303), .O(\uart_tx_inst/n858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6454.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6455 (.I0(n2326), .I1(\uart_tx_inst/r_Clock_Count [24]), 
            .I2(\uart_tx_inst/r_Clock_Count [25]), .O(n2328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6455.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6456 (.I0(n2325), .I1(n2328), .I2(\uart_tx_inst/r_Clock_Count [26]), 
            .I3(n2303), .O(\uart_tx_inst/n861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6456.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6457 (.I0(n2324), .I1(n2328), .I2(\uart_tx_inst/r_Clock_Count [26]), 
            .O(n2329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6457.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6458 (.I0(n2321), .I1(n2329), .I2(\uart_tx_inst/r_Clock_Count [27]), 
            .I3(n2303), .O(\uart_tx_inst/n864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6458.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6459 (.I0(n2324), .I1(n2328), .I2(\uart_tx_inst/r_Clock_Count [26]), 
            .I3(\uart_tx_inst/r_Clock_Count [27]), .O(n2330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6459.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6460 (.I0(n2318), .I1(n2330), .I2(n2320), .O(n2331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6460.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6461 (.I0(n2331), .I1(\uart_tx_inst/r_Clock_Count [28]), 
            .I2(n2303), .O(\uart_tx_inst/n867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6461.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6462 (.I0(n2331), .I1(\uart_tx_inst/r_Clock_Count [28]), 
            .I2(\uart_tx_inst/r_Clock_Count [29]), .I3(n2303), .O(\uart_tx_inst/n870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6462.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6463 (.I0(\uart_tx_inst/r_Clock_Count [28]), .I1(\uart_tx_inst/r_Clock_Count [29]), 
            .O(n2332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6463.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6464 (.I0(n2331), .I1(n2332), .I2(\uart_tx_inst/r_Clock_Count [30]), 
            .I3(n2303), .O(\uart_tx_inst/n873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6464.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6465 (.I0(n2332), .I1(\uart_tx_inst/r_Clock_Count [12]), 
            .I2(\uart_tx_inst/r_Clock_Count [13]), .I3(\uart_tx_inst/r_Clock_Count [30]), 
            .O(n2333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6465.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6466 (.I0(n2333), .I1(n2320), .O(n2334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6466.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6467 (.I0(n2313), .I1(n2330), .I2(n2334), .I3(n2315), 
            .O(n2335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6467.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6468 (.I0(n2335), .I1(\uart_tx_inst/r_Clock_Count [31]), 
            .I2(n2303), .O(\uart_tx_inst/n876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(240)
    defparam LUT__6468.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6469 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_SM_Main [1]), .O(\uart_tx_inst/n880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(260)
    defparam LUT__6469.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6470 (.I0(\uart_tx_inst/r_Bit_Index [0]), .I1(\uart_tx_inst/r_Bit_Index [1]), 
            .I2(\uart_tx_inst/r_Bit_Index [2]), .I3(\uart_tx_inst/r_SM_Main [1]), 
            .O(\uart_tx_inst/n884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(260)
    defparam LUT__6470.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6471 (.I0(\uart_tx_inst/r_SM_Main [2]), .I1(n2292), .O(\uart_tx_inst/n1032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(44)
    defparam LUT__6471.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__6472 (.I0(\uart_tx_inst/r_SM_Main [0]), .I1(\uart_tx_inst/r_SM_Main [2]), 
            .I2(n2309), .O(\uart_tx_inst/n1224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(44)
    defparam LUT__6472.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6473 (.I0(\uart_tx_inst/n50 ), .I1(\uart_tx_inst/r_SM_Main [0]), 
            .I2(\uart_tx_inst/r_SM_Main [1]), .O(\uart_tx_inst/n779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(287)
    defparam LUT__6473.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__6474 (.I0(\uart_tx_inst/r_SM_Main [2]), .I1(\uart_tx_inst/r_SM_Main [1]), 
            .I2(\uart_tx_inst/r_SM_Main [0]), .O(\uart_tx_inst/n1206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(44)
    defparam LUT__6474.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6475 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [5]), 
            .O(rx_data[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6475.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6476 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [6]), 
            .O(rx_data[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6476.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6477 (.I0(rx_ready), .I1(\uart_rx_inst/r_Rx_Byte [7]), 
            .O(rx_data[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6477.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6480 (.I0(tx_2), .O(tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(288)
    defparam LUT__6480.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__6229 (.I0(\uart_rx_inst/r_Rx_Byte [0]), .I1(rx_ready), 
            .O(rx_data[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/half_adder.v(171)
    defparam LUT__6229.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter [0]), 
            .I1(1'b1), .CI(1'b0), .CO(n2337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4646)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt [0]), 
            .I1(1'b1), .CI(1'b0), .CO(n2336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/trinity/Downloads/efinity/2024.2/project/verilog_learnings/work_dbg/debug_top.v(4660)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_bbdc1861_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_bbdc1861_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bbdc1861__5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_bbdc1861__5_5_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_bbdc1861_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_bbdc1861_0
// module not written out since it is a black box. 
//

