module add_gate(
input a, b,
output sum
);

assign sum= a + b;

endmodule
